module ALU(
  input  [3:0]  io_fn,
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_alu_out,
  output        io_cmp_out
);
  wire [31:0] _in2_inv_T_1 = ~io_in2; // @[ALU.scala 90:35]
  wire [31:0] in2_inv = io_fn[3] ? _in2_inv_T_1 : io_in2; // @[ALU.scala 90:20]
  wire [31:0] in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 92:28]
  wire [31:0] _adder_out_T_1 = io_in1 + in2_inv; // @[ALU.scala 93:26]
  wire [31:0] _GEN_0 = {{31'd0}, io_fn[3]}; // @[ALU.scala 93:36]
  wire [31:0] adder_out = _adder_out_T_1 + _GEN_0; // @[ALU.scala 93:36]
  wire  _slt_T_2 = io_in1[31] == io_in2[31]; // @[ALU.scala 98:18]
  wire  _slt_T_7 = io_fn[1] ? io_in2[31] : io_in1[31]; // @[ALU.scala 100:10]
  wire  slt = _slt_T_2 ? adder_out[31] : _slt_T_7; // @[ALU.scala 97:8]
  wire  _io_cmp_out_T_2 = ~io_fn[3]; // @[ALU.scala 66:26]
  wire  _io_cmp_out_T_4 = _io_cmp_out_T_2 ? in1_xor_in2 == 32'h0 : slt; // @[ALU.scala 102:41]
  wire [4:0] shamt = io_in2[4:0]; // @[ALU.scala 105:32]
  wire  _shin_T_2 = io_fn == 4'h5 | io_fn == 4'hb; // @[ALU.scala 106:34]
  wire [31:0] _GEN_1 = {{16'd0}, io_in1[31:16]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_6 = _GEN_1 & 32'hffff; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_8 = {io_in1[15:0], 16'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_10 = _shin_T_8 & 32'hffff0000; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_11 = _shin_T_6 | _shin_T_10; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_2 = {{8'd0}, _shin_T_11[31:8]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_16 = _GEN_2 & 32'hff00ff; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_18 = {_shin_T_11[23:0], 8'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_20 = _shin_T_18 & 32'hff00ff00; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_21 = _shin_T_16 | _shin_T_20; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_3 = {{4'd0}, _shin_T_21[31:4]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_26 = _GEN_3 & 32'hf0f0f0f; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_28 = {_shin_T_21[27:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_30 = _shin_T_28 & 32'hf0f0f0f0; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_31 = _shin_T_26 | _shin_T_30; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_4 = {{2'd0}, _shin_T_31[31:2]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_36 = _GEN_4 & 32'h33333333; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_38 = {_shin_T_31[29:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_40 = _shin_T_38 & 32'hcccccccc; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_41 = _shin_T_36 | _shin_T_40; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_5 = {{1'd0}, _shin_T_41[31:1]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_46 = _GEN_5 & 32'h55555555; // @[Bitwise.scala 105:31]
  wire [31:0] _shin_T_48 = {_shin_T_41[30:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shin_T_50 = _shin_T_48 & 32'haaaaaaaa; // @[Bitwise.scala 105:80]
  wire [31:0] _shin_T_51 = _shin_T_46 | _shin_T_50; // @[Bitwise.scala 105:39]
  wire [31:0] shin = io_fn == 4'h5 | io_fn == 4'hb ? io_in1 : _shin_T_51; // @[ALU.scala 106:17]
  wire  _shout_r_T_2 = io_fn[3] & shin[31]; // @[ALU.scala 107:35]
  wire [32:0] _shout_r_T_4 = {_shout_r_T_2,shin}; // @[ALU.scala 107:53]
  wire [32:0] _shout_r_T_5 = $signed(_shout_r_T_4) >>> shamt; // @[ALU.scala 107:60]
  wire [31:0] shout_r = _shout_r_T_5[31:0]; // @[ALU.scala 107:69]
  wire [31:0] _GEN_6 = {{16'd0}, shout_r[31:16]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_3 = _GEN_6 & 32'hffff; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_5 = {shout_r[15:0], 16'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_7 = _shout_l_T_5 & 32'hffff0000; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_8 = _shout_l_T_3 | _shout_l_T_7; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_7 = {{8'd0}, _shout_l_T_8[31:8]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_13 = _GEN_7 & 32'hff00ff; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_15 = {_shout_l_T_8[23:0], 8'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_17 = _shout_l_T_15 & 32'hff00ff00; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_18 = _shout_l_T_13 | _shout_l_T_17; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_8 = {{4'd0}, _shout_l_T_18[31:4]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_23 = _GEN_8 & 32'hf0f0f0f; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_25 = {_shout_l_T_18[27:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_27 = _shout_l_T_25 & 32'hf0f0f0f0; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_28 = _shout_l_T_23 | _shout_l_T_27; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_9 = {{2'd0}, _shout_l_T_28[31:2]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_33 = _GEN_9 & 32'h33333333; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_35 = {_shout_l_T_28[29:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_37 = _shout_l_T_35 & 32'hcccccccc; // @[Bitwise.scala 105:80]
  wire [31:0] _shout_l_T_38 = _shout_l_T_33 | _shout_l_T_37; // @[Bitwise.scala 105:39]
  wire [31:0] _GEN_10 = {{1'd0}, _shout_l_T_38[31:1]}; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_43 = _GEN_10 & 32'h55555555; // @[Bitwise.scala 105:31]
  wire [31:0] _shout_l_T_45 = {_shout_l_T_38[30:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [31:0] _shout_l_T_47 = _shout_l_T_45 & 32'haaaaaaaa; // @[Bitwise.scala 105:80]
  wire [31:0] shout_l = _shout_l_T_43 | _shout_l_T_47; // @[Bitwise.scala 105:39]
  wire [31:0] _shout_T_3 = _shin_T_2 ? shout_r : 32'h0; // @[ALU.scala 109:18]
  wire [31:0] _shout_T_5 = io_fn == 4'h1 ? shout_l : 32'h0; // @[ALU.scala 110:8]
  wire [31:0] shout = _shout_T_3 | _shout_T_5; // @[ALU.scala 109:70]
  wire  _logic_T_1 = io_fn == 4'h6; // @[ALU.scala 113:45]
  wire [31:0] _logic_T_3 = io_fn == 4'h4 | io_fn == 4'h6 ? in1_xor_in2 : 32'h0; // @[ALU.scala 113:18]
  wire [31:0] _logic_T_7 = io_in1 & io_in2; // @[ALU.scala 114:53]
  wire [31:0] _logic_T_8 = _logic_T_1 | io_fn == 4'h7 ? _logic_T_7 : 32'h0; // @[ALU.scala 114:8]
  wire [31:0] logic_ = _logic_T_3 | _logic_T_8; // @[ALU.scala 113:74]
  wire  _shift_logic_T = io_fn >= 4'hc; // @[ALU.scala 52:30]
  wire  _shift_logic_T_1 = _shift_logic_T & slt; // @[ALU.scala 115:35]
  wire [31:0] _GEN_11 = {{31'd0}, _shift_logic_T_1}; // @[ALU.scala 115:43]
  wire [31:0] _shift_logic_T_2 = _GEN_11 | logic_; // @[ALU.scala 115:43]
  wire [31:0] shift_logic = _shift_logic_T_2 | shout; // @[ALU.scala 115:51]
  assign io_alu_out = io_fn == 4'h0 | io_fn == 4'ha ? adder_out : shift_logic; // @[ALU.scala 117:8]
  assign io_cmp_out = io_fn[0] ^ _io_cmp_out_T_4; // @[ALU.scala 102:36]
endmodule
module RISCV(
  input         clock,
  input         reset,
  output [31:0] io_iData_addr,
  input  [31:0] io_iData_inst,
  output [31:0] io_dData_addr,
  output [31:0] io_dData_writeData,
  output        io_dData_writeEnable,
  input  [31:0] io_dData_readData
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] rf [0:31]; // @[Register.scala 8:15]
  wire  rf_id_rs_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_id_rs_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_id_rs_MPORT_data; // @[Register.scala 8:15]
  wire  rf_id_rs_MPORT_1_en; // @[Register.scala 8:15]
  wire [4:0] rf_id_rs_MPORT_1_addr; // @[Register.scala 8:15]
  wire [31:0] rf_id_rs_MPORT_1_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_0_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_0_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_0_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_1_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_1_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_1_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_2_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_2_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_2_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_3_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_3_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_3_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_4_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_4_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_4_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_5_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_5_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_5_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_6_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_6_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_6_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_7_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_7_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_7_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_8_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_8_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_8_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_9_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_9_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_9_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_10_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_10_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_10_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_11_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_11_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_11_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_12_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_12_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_12_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_13_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_13_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_13_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_14_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_14_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_14_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_15_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_15_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_15_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_16_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_16_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_16_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_17_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_17_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_17_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_18_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_18_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_18_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_19_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_19_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_19_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_20_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_20_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_20_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_21_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_21_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_21_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_22_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_22_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_22_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_23_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_23_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_23_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_24_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_24_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_24_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_25_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_25_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_25_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_26_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_26_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_26_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_27_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_27_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_27_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_28_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_28_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_28_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_29_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_29_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_29_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_30_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_30_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_30_MPORT_data; // @[Register.scala 8:15]
  wire  rf_io_dbg_monitor_reg_31_MPORT_en; // @[Register.scala 8:15]
  wire [4:0] rf_io_dbg_monitor_reg_31_MPORT_addr; // @[Register.scala 8:15]
  wire [31:0] rf_io_dbg_monitor_reg_31_MPORT_data; // @[Register.scala 8:15]
  wire [31:0] rf_MPORT_data; // @[Register.scala 8:15]
  wire [4:0] rf_MPORT_addr; // @[Register.scala 8:15]
  wire  rf_MPORT_mask; // @[Register.scala 8:15]
  wire  rf_MPORT_en; // @[Register.scala 8:15]
  wire  rf_clock;
  wire [3:0] alu_io_fn; // @[RISCV.scala 289:19]
  wire [31:0] alu_io_in1; // @[RISCV.scala 289:19]
  wire [31:0] alu_io_in2; // @[RISCV.scala 289:19]
  wire [31:0] alu_io_alu_out; // @[RISCV.scala 289:19]
  wire  alu_io_cmp_out; // @[RISCV.scala 289:19]
  reg [31:0] id_pc; // @[RISCV.scala 58:22]
  reg [31:0] id_npc; // @[RISCV.scala 59:23]
  reg [31:0] id_inst; // @[RISCV.scala 60:24]
  reg [31:0] ex_pc; // @[RISCV.scala 70:22]
  reg [31:0] ex_npc; // @[RISCV.scala 71:23]
  reg [31:0] ex_inst; // @[RISCV.scala 72:24]
  reg  ex_ctrl_branch; // @[RISCV.scala 73:24]
  reg  ex_ctrl_jal; // @[RISCV.scala 73:24]
  reg  ex_ctrl_jalr; // @[RISCV.scala 73:24]
  reg [1:0] ex_ctrl_sel_alu1; // @[RISCV.scala 73:24]
  reg [1:0] ex_ctrl_sel_alu2; // @[RISCV.scala 73:24]
  reg [2:0] ex_ctrl_sel_imm; // @[RISCV.scala 73:24]
  reg [3:0] ex_ctrl_alu_fn; // @[RISCV.scala 73:24]
  reg  ex_ctrl_mem; // @[RISCV.scala 73:24]
  reg [4:0] ex_ctrl_mem_cmd; // @[RISCV.scala 73:24]
  reg  ex_ctrl_wxd; // @[RISCV.scala 73:24]
  reg [4:0] ex_reg_raddr_0; // @[RISCV.scala 74:29]
  reg [4:0] ex_reg_raddr_1; // @[RISCV.scala 74:29]
  reg [4:0] ex_reg_waddr; // @[RISCV.scala 75:29]
  reg [31:0] ex_rs_0; // @[RISCV.scala 76:22]
  reg [31:0] ex_rs_1; // @[RISCV.scala 76:22]
  reg [31:0] mem_pc; // @[RISCV.scala 87:23]
  reg [31:0] mem_npc; // @[RISCV.scala 88:24]
  reg  mem_ctrl_branch; // @[RISCV.scala 89:25]
  reg  mem_ctrl_jal; // @[RISCV.scala 89:25]
  reg  mem_ctrl_jalr; // @[RISCV.scala 89:25]
  reg  mem_ctrl_mem; // @[RISCV.scala 89:25]
  reg [4:0] mem_ctrl_mem_cmd; // @[RISCV.scala 89:25]
  reg  mem_ctrl_wxd; // @[RISCV.scala 89:25]
  reg [4:0] mem_reg_waddr; // @[RISCV.scala 90:30]
  reg [31:0] mem_rs_1; // @[RISCV.scala 91:23]
  reg [31:0] mem_imm; // @[RISCV.scala 92:24]
  reg [31:0] mem_alu_out; // @[RISCV.scala 93:28]
  reg  mem_alu_cmp_out; // @[RISCV.scala 94:32]
  reg [31:0] wb_npc; // @[RISCV.scala 102:23]
  reg  wb_ctrl_jalr; // @[RISCV.scala 103:24]
  reg  wb_ctrl_mem; // @[RISCV.scala 103:24]
  reg  wb_ctrl_wxd; // @[RISCV.scala 103:24]
  reg [4:0] wb_reg_waddr; // @[RISCV.scala 105:29]
  reg [31:0] wb_alu_out; // @[RISCV.scala 106:27]
  reg [31:0] wb_dData_readData; // @[RISCV.scala 107:34]
  reg [31:0] pc; // @[RISCV.scala 127:19]
  wire [31:0] npc = pc + 32'h4; // @[RISCV.scala 131:13]
  wire [4:0] id_inst_arange_rs1 = id_inst[19:15]; // @[Decode.scala 19:20]
  wire [4:0] id_inst_arange_rs2 = id_inst[24:20]; // @[Decode.scala 20:20]
  wire  _load_stall_T_2 = id_inst_arange_rs1 == ex_reg_waddr | id_inst_arange_rs2 == ex_reg_waddr; // @[RISCV.scala 192:48]
  wire  load_stall = _load_stall_T_2 & ex_ctrl_mem & ex_ctrl_mem_cmd == 5'h0; // @[RISCV.scala 193:28]
  wire  _T = ~load_stall; // @[RISCV.scala 152:8]
  wire  _jump_flush_T_5 = mem_ctrl_branch & mem_alu_cmp_out | mem_ctrl_jal; // @[RISCV.scala 342:63]
  wire  jump_flush = mem_ctrl_branch & mem_alu_cmp_out | mem_ctrl_jal | mem_ctrl_jalr; // @[RISCV.scala 342:87]
  wire  _T_1 = ~jump_flush; // @[RISCV.scala 152:23]
  wire  _T_2 = ~load_stall & ~jump_flush; // @[RISCV.scala 152:20]
  wire [4:0] id_inst_arange_rd = id_inst[11:7]; // @[Decode.scala 18:19]
  wire [31:0] _id_ctrl_decoder_ctrl_signals_T = id_inst & 32'h707f; // @[RetentionBundle.scala 170:15]
  wire  id_ctrl_decoder_0 = 32'h63 == _id_ctrl_decoder_ctrl_signals_T; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_3 = 32'h67 == _id_ctrl_decoder_ctrl_signals_T; // @[RetentionBundle.scala 170:15]
  wire [31:0] _id_ctrl_decoder_ctrl_signals_T_4 = id_inst & 32'h7f; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_5 = 32'h6f == _id_ctrl_decoder_ctrl_signals_T_4; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_7 = 32'h37 == _id_ctrl_decoder_ctrl_signals_T_4; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_9 = 32'h17 == _id_ctrl_decoder_ctrl_signals_T_4; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_11 = 32'h13 == _id_ctrl_decoder_ctrl_signals_T; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_13 = 32'h3 == _id_ctrl_decoder_ctrl_signals_T; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_15 = 32'h23 == _id_ctrl_decoder_ctrl_signals_T; // @[RetentionBundle.scala 170:15]
  wire  _id_ctrl_decoder_ctrl_signals_T_45 = _id_ctrl_decoder_ctrl_signals_T_3 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_5; // @[Mux.scala 101:16]
  wire  id_ctrl_decoder_1 = id_ctrl_decoder_0 ? 1'h0 : _id_ctrl_decoder_ctrl_signals_T_45; // @[Mux.scala 101:16]
  wire  id_ctrl_decoder_2 = id_ctrl_decoder_0 ? 1'h0 : _id_ctrl_decoder_ctrl_signals_T_3; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_87 = _id_ctrl_decoder_ctrl_signals_T_11 | (_id_ctrl_decoder_ctrl_signals_T_13 |
    _id_ctrl_decoder_ctrl_signals_T_15); // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_88 = _id_ctrl_decoder_ctrl_signals_T_9 ? 2'h2 : {{1'd0},
    _id_ctrl_decoder_ctrl_signals_T_87}; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_89 = _id_ctrl_decoder_ctrl_signals_T_7 ? 2'h0 :
    _id_ctrl_decoder_ctrl_signals_T_88; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_90 = _id_ctrl_decoder_ctrl_signals_T_5 ? 2'h2 :
    _id_ctrl_decoder_ctrl_signals_T_89; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_108 = _id_ctrl_decoder_ctrl_signals_T_15 ? 2'h3 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_109 = _id_ctrl_decoder_ctrl_signals_T_13 ? 2'h3 :
    _id_ctrl_decoder_ctrl_signals_T_108; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_110 = _id_ctrl_decoder_ctrl_signals_T_11 ? 2'h3 :
    _id_ctrl_decoder_ctrl_signals_T_109; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_111 = _id_ctrl_decoder_ctrl_signals_T_9 ? 2'h3 :
    _id_ctrl_decoder_ctrl_signals_T_110; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_112 = _id_ctrl_decoder_ctrl_signals_T_7 ? 2'h3 :
    _id_ctrl_decoder_ctrl_signals_T_111; // @[Mux.scala 101:16]
  wire [1:0] _id_ctrl_decoder_ctrl_signals_T_113 = _id_ctrl_decoder_ctrl_signals_T_5 ? 2'h1 :
    _id_ctrl_decoder_ctrl_signals_T_112; // @[Mux.scala 101:16]
  wire [2:0] _id_ctrl_decoder_ctrl_signals_T_132 = _id_ctrl_decoder_ctrl_signals_T_13 ? 3'h4 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _id_ctrl_decoder_ctrl_signals_T_133 = _id_ctrl_decoder_ctrl_signals_T_11 ? 3'h4 :
    _id_ctrl_decoder_ctrl_signals_T_132; // @[Mux.scala 101:16]
  wire [2:0] _id_ctrl_decoder_ctrl_signals_T_134 = _id_ctrl_decoder_ctrl_signals_T_9 ? 3'h2 :
    _id_ctrl_decoder_ctrl_signals_T_133; // @[Mux.scala 101:16]
  wire [2:0] _id_ctrl_decoder_ctrl_signals_T_135 = _id_ctrl_decoder_ctrl_signals_T_7 ? 3'h2 :
    _id_ctrl_decoder_ctrl_signals_T_134; // @[Mux.scala 101:16]
  wire [2:0] _id_ctrl_decoder_ctrl_signals_T_136 = _id_ctrl_decoder_ctrl_signals_T_5 ? 3'h3 :
    _id_ctrl_decoder_ctrl_signals_T_135; // @[Mux.scala 101:16]
  wire [1:0] id_ctrl_decoder_6 = id_ctrl_decoder_0 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_179 = _id_ctrl_decoder_ctrl_signals_T_11 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_13 | _id_ctrl_decoder_ctrl_signals_T_15; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_180 = _id_ctrl_decoder_ctrl_signals_T_9 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_179; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_181 = _id_ctrl_decoder_ctrl_signals_T_7 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_180; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_182 = _id_ctrl_decoder_ctrl_signals_T_5 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_181; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_183 = _id_ctrl_decoder_ctrl_signals_T_3 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_182; // @[Mux.scala 101:16]
  wire  id_ctrl_decoder_7 = id_ctrl_decoder_0 ? 1'h0 : _id_ctrl_decoder_ctrl_signals_T_183; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_201 = _id_ctrl_decoder_ctrl_signals_T_13 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_15; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_202 = _id_ctrl_decoder_ctrl_signals_T_11 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_201; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_203 = _id_ctrl_decoder_ctrl_signals_T_9 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_202; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_204 = _id_ctrl_decoder_ctrl_signals_T_7 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_203; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_205 = _id_ctrl_decoder_ctrl_signals_T_5 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_204; // @[Mux.scala 101:16]
  wire  _id_ctrl_decoder_ctrl_signals_T_206 = _id_ctrl_decoder_ctrl_signals_T_3 ? 1'h0 :
    _id_ctrl_decoder_ctrl_signals_T_205; // @[Mux.scala 101:16]
  wire  id_ctrl_decoder_8 = id_ctrl_decoder_0 ? 1'h0 : _id_ctrl_decoder_ctrl_signals_T_206; // @[Mux.scala 101:16]
  wire  id_ctrl_decoder_10 = id_ctrl_decoder_0 ? 1'h0 : _id_ctrl_decoder_ctrl_signals_T_3 | (
    _id_ctrl_decoder_ctrl_signals_T_5 | (_id_ctrl_decoder_ctrl_signals_T_7 | (_id_ctrl_decoder_ctrl_signals_T_9 | (
    _id_ctrl_decoder_ctrl_signals_T_11 | _id_ctrl_decoder_ctrl_signals_T_13)))); // @[Mux.scala 101:16]
  wire  _GEN_9 = _T_2 ? id_ctrl_decoder_10 : 1'h1; // @[RISCV.scala 212:36 216:13 223:13]
  wire [4:0] id_ctrl_mem_cmd = {{4'd0}, id_ctrl_decoder_8}; // @[RISCV.scala 172:9 RetentionBundle.scala 90:56]
  wire  _GEN_12 = _T_2 & id_ctrl_decoder_7; // @[RISCV.scala 212:36 216:13 223:13]
  wire [3:0] id_ctrl_alu_fn = {{2'd0}, id_ctrl_decoder_6}; // @[RISCV.scala 172:9 RetentionBundle.scala 90:56]
  wire  _GEN_17 = _T_2 & id_ctrl_decoder_2; // @[RISCV.scala 212:36 216:13 223:13]
  wire  _GEN_18 = _T_2 & id_ctrl_decoder_1; // @[RISCV.scala 212:36 216:13 223:13]
  wire  _GEN_19 = _T_2 & id_ctrl_decoder_0; // @[RISCV.scala 212:36 216:13 223:13]
  wire  _ex_rs_bypassed_T = ex_reg_raddr_0 != 5'h0; // @[RISCV.scala 240:29]
  wire  _ex_rs_bypassed_T_2 = _ex_rs_bypassed_T & ex_reg_raddr_0 == mem_reg_waddr; // @[RISCV.scala 241:13]
  wire  _ex_rs_bypassed_T_5 = _ex_rs_bypassed_T_2 & mem_ctrl_wxd; // @[RISCV.scala 242:13]
  wire  _ex_rs_bypassed_T_8 = _ex_rs_bypassed_T & ex_reg_raddr_0 == wb_reg_waddr; // @[RISCV.scala 247:13]
  wire  _ex_rs_bypassed_T_11 = _ex_rs_bypassed_T_8 & wb_ctrl_wxd; // @[RISCV.scala 248:13]
  wire  _ex_rs_bypassed_T_14 = _ex_rs_bypassed_T_11 & wb_ctrl_mem; // @[RISCV.scala 249:13]
  wire [31:0] _ex_rs_bypassed_T_15 = _ex_rs_bypassed_T_14 ? io_dData_readData : ex_rs_0; // @[Mux.scala 101:16]
  wire [31:0] ex_rs_bypassed_0 = _ex_rs_bypassed_T_5 ? mem_alu_out : _ex_rs_bypassed_T_15; // @[Mux.scala 101:16]
  wire  _ex_rs_bypassed_T_16 = ex_reg_raddr_1 != 5'h0; // @[RISCV.scala 240:29]
  wire  _ex_rs_bypassed_T_18 = _ex_rs_bypassed_T_16 & ex_reg_raddr_1 == mem_reg_waddr; // @[RISCV.scala 241:13]
  wire  _ex_rs_bypassed_T_21 = _ex_rs_bypassed_T_18 & mem_ctrl_wxd; // @[RISCV.scala 242:13]
  wire  _ex_rs_bypassed_T_24 = _ex_rs_bypassed_T_16 & ex_reg_raddr_1 == wb_reg_waddr; // @[RISCV.scala 247:13]
  wire  _ex_rs_bypassed_T_27 = _ex_rs_bypassed_T_24 & wb_ctrl_wxd; // @[RISCV.scala 248:13]
  wire  _ex_rs_bypassed_T_30 = _ex_rs_bypassed_T_27 & wb_ctrl_mem; // @[RISCV.scala 249:13]
  wire [31:0] _ex_rs_bypassed_T_31 = _ex_rs_bypassed_T_30 ? io_dData_readData : ex_rs_1; // @[Mux.scala 101:16]
  wire [31:0] ex_rs_bypassed_1 = _ex_rs_bypassed_T_21 ? mem_alu_out : _ex_rs_bypassed_T_31; // @[Mux.scala 101:16]
  wire  _ex_imm_sign_T = ex_ctrl_sel_imm == 3'h5; // @[ImmGenerate.scala 20:24]
  wire  _ex_imm_sign_T_2 = ex_inst[31]; // @[ImmGenerate.scala 20:49]
  wire  ex_imm_sign = ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2); // @[ImmGenerate.scala 20:19]
  wire  _ex_imm_b30_20_T = ex_ctrl_sel_imm == 3'h2; // @[ImmGenerate.scala 21:26]
  wire [10:0] _ex_imm_b30_20_T_2 = ex_inst[30:20]; // @[ImmGenerate.scala 21:50]
  wire [7:0] _ex_imm_b19_12_T_4 = ex_inst[19:12]; // @[ImmGenerate.scala 22:73]
  wire  _ex_imm_b11_T_2 = _ex_imm_b30_20_T | _ex_imm_sign_T; // @[ImmGenerate.scala 24:21]
  wire  _ex_imm_b11_T_3 = ex_ctrl_sel_imm == 3'h3; // @[ImmGenerate.scala 27:13]
  wire  _ex_imm_b11_T_5 = ex_inst[20]; // @[ImmGenerate.scala 28:18]
  wire  _ex_imm_b11_T_6 = ex_ctrl_sel_imm == 3'h1; // @[ImmGenerate.scala 29:17]
  wire  _ex_imm_b11_T_8 = ex_inst[7]; // @[ImmGenerate.scala 29:36]
  wire  _ex_imm_b11_T_9 = ex_ctrl_sel_imm == 3'h1 ? $signed(_ex_imm_b11_T_8) : $signed(ex_imm_sign); // @[ImmGenerate.scala 29:12]
  wire  _ex_imm_b11_T_10 = _ex_imm_b11_T_3 ? $signed(_ex_imm_b11_T_5) : $signed(_ex_imm_b11_T_9); // @[ImmGenerate.scala 26:10]
  wire [5:0] ex_imm_b10_5 = _ex_imm_b11_T_2 ? 6'h0 : ex_inst[30:25]; // @[ImmGenerate.scala 32:20]
  wire  _ex_imm_b4_1_T_1 = ex_ctrl_sel_imm == 3'h0; // @[ImmGenerate.scala 37:13]
  wire  _ex_imm_b4_1_T_3 = ex_ctrl_sel_imm == 3'h0 | _ex_imm_b11_T_6; // @[ImmGenerate.scala 37:23]
  wire [3:0] _ex_imm_b4_1_T_8 = _ex_imm_sign_T ? ex_inst[19:16] : ex_inst[24:21]; // @[ImmGenerate.scala 39:12]
  wire [3:0] _ex_imm_b4_1_T_9 = _ex_imm_b4_1_T_3 ? ex_inst[11:8] : _ex_imm_b4_1_T_8; // @[ImmGenerate.scala 36:10]
  wire [3:0] ex_imm_b4_1 = _ex_imm_b30_20_T ? 4'h0 : _ex_imm_b4_1_T_9; // @[ImmGenerate.scala 33:19]
  wire  _ex_imm_b0_T_7 = ex_ctrl_sel_imm == 3'h4 ? ex_inst[20] : _ex_imm_sign_T & ex_inst[15]; // @[ImmGenerate.scala 45:10]
  wire  ex_imm_b0 = _ex_imm_b4_1_T_1 ? ex_inst[7] : _ex_imm_b0_T_7; // @[ImmGenerate.scala 42:17]
  wire  ex_imm_hi_lo_lo = _ex_imm_b11_T_2 ? $signed(1'sh0) : $signed(_ex_imm_b11_T_10); // @[Cat.scala 31:58]
  wire [7:0] ex_imm_hi_lo_hi = ex_ctrl_sel_imm != 3'h2 & ex_ctrl_sel_imm != 3'h3 ? $signed({8{ex_imm_sign}}) : $signed(
    _ex_imm_b19_12_T_4); // @[Cat.scala 31:58]
  wire [10:0] ex_imm_hi_hi_lo = ex_ctrl_sel_imm == 3'h2 ? $signed(_ex_imm_b30_20_T_2) : $signed({11{ex_imm_sign}}); // @[Cat.scala 31:58]
  wire  ex_imm_hi_hi_hi = ex_ctrl_sel_imm == 3'h5 ? $signed(1'sh0) : $signed(_ex_imm_sign_T_2); // @[Cat.scala 31:58]
  wire [31:0] ex_imm = {ex_imm_hi_hi_hi,ex_imm_hi_hi_lo,ex_imm_hi_lo_hi,ex_imm_hi_lo_lo,ex_imm_b10_5,ex_imm_b4_1,
    ex_imm_b0}; // @[ImmGenerate.scala 48:53]
  wire [31:0] _ex_op1_T_1 = 2'h1 == ex_ctrl_sel_alu1 ? ex_rs_bypassed_0 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _ex_op2_T = {ex_imm_hi_hi_hi,ex_imm_hi_hi_lo,ex_imm_hi_lo_hi,ex_imm_hi_lo_lo,ex_imm_b10_5,ex_imm_b4_1,
    ex_imm_b0}; // @[RISCV.scala 281:25]
  wire [31:0] _ex_op2_T_2 = 2'h2 == ex_ctrl_sel_alu2 ? ex_rs_bypassed_1 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _ex_op2_T_4 = 2'h3 == ex_ctrl_sel_alu2 ? _ex_op2_T : _ex_op2_T_2; // @[Mux.scala 81:58]
  wire  _GEN_27 = _T_1 ? ex_ctrl_wxd : 1'h1; // @[RISCV.scala 308:21 311:14 320:14]
  wire  _GEN_30 = _T_1 & ex_ctrl_mem; // @[RISCV.scala 308:21 311:14 320:14]
  wire  _GEN_35 = _T_1 & ex_ctrl_jalr; // @[RISCV.scala 308:21 311:14 320:14]
  wire  _GEN_36 = _T_1 & ex_ctrl_jal; // @[RISCV.scala 308:21 311:14 320:14]
  wire  _GEN_37 = _T_1 & ex_ctrl_branch; // @[RISCV.scala 308:21 311:14 320:14]
  wire  _GEN_43 = _T_1 & alu_io_cmp_out; // @[RISCV.scala 308:21 316:21 325:21]
  wire [31:0] _rf_wdata_T_4 = wb_ctrl_mem ? wb_dData_readData : wb_alu_out; // @[Mux.scala 101:16]
  wire  _T_7 = wb_reg_waddr != 5'h0; // @[Register.scala 17:15]
  wire [31:0] _pc_T_8 = mem_pc + mem_imm; // @[RISCV.scala 387:89]
  ALU alu ( // @[RISCV.scala 289:19]
    .io_fn(alu_io_fn),
    .io_in1(alu_io_in1),
    .io_in2(alu_io_in2),
    .io_alu_out(alu_io_alu_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  assign rf_id_rs_MPORT_en = 1'h1;
  assign rf_id_rs_MPORT_addr = id_inst[19:15];
  assign rf_id_rs_MPORT_data = rf[rf_id_rs_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_id_rs_MPORT_1_en = 1'h1;
  assign rf_id_rs_MPORT_1_addr = id_inst[24:20];
  assign rf_id_rs_MPORT_1_data = rf[rf_id_rs_MPORT_1_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_0_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_0_MPORT_addr = 5'h0;
  assign rf_io_dbg_monitor_reg_0_MPORT_data = rf[rf_io_dbg_monitor_reg_0_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_1_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_1_MPORT_addr = 5'h1;
  assign rf_io_dbg_monitor_reg_1_MPORT_data = rf[rf_io_dbg_monitor_reg_1_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_2_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_2_MPORT_addr = 5'h2;
  assign rf_io_dbg_monitor_reg_2_MPORT_data = rf[rf_io_dbg_monitor_reg_2_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_3_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_3_MPORT_addr = 5'h3;
  assign rf_io_dbg_monitor_reg_3_MPORT_data = rf[rf_io_dbg_monitor_reg_3_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_4_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_4_MPORT_addr = 5'h4;
  assign rf_io_dbg_monitor_reg_4_MPORT_data = rf[rf_io_dbg_monitor_reg_4_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_5_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_5_MPORT_addr = 5'h5;
  assign rf_io_dbg_monitor_reg_5_MPORT_data = rf[rf_io_dbg_monitor_reg_5_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_6_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_6_MPORT_addr = 5'h6;
  assign rf_io_dbg_monitor_reg_6_MPORT_data = rf[rf_io_dbg_monitor_reg_6_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_7_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_7_MPORT_addr = 5'h7;
  assign rf_io_dbg_monitor_reg_7_MPORT_data = rf[rf_io_dbg_monitor_reg_7_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_8_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_8_MPORT_addr = 5'h8;
  assign rf_io_dbg_monitor_reg_8_MPORT_data = rf[rf_io_dbg_monitor_reg_8_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_9_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_9_MPORT_addr = 5'h9;
  assign rf_io_dbg_monitor_reg_9_MPORT_data = rf[rf_io_dbg_monitor_reg_9_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_10_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_10_MPORT_addr = 5'ha;
  assign rf_io_dbg_monitor_reg_10_MPORT_data = rf[rf_io_dbg_monitor_reg_10_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_11_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_11_MPORT_addr = 5'hb;
  assign rf_io_dbg_monitor_reg_11_MPORT_data = rf[rf_io_dbg_monitor_reg_11_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_12_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_12_MPORT_addr = 5'hc;
  assign rf_io_dbg_monitor_reg_12_MPORT_data = rf[rf_io_dbg_monitor_reg_12_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_13_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_13_MPORT_addr = 5'hd;
  assign rf_io_dbg_monitor_reg_13_MPORT_data = rf[rf_io_dbg_monitor_reg_13_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_14_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_14_MPORT_addr = 5'he;
  assign rf_io_dbg_monitor_reg_14_MPORT_data = rf[rf_io_dbg_monitor_reg_14_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_15_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_15_MPORT_addr = 5'hf;
  assign rf_io_dbg_monitor_reg_15_MPORT_data = rf[rf_io_dbg_monitor_reg_15_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_16_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_16_MPORT_addr = 5'h10;
  assign rf_io_dbg_monitor_reg_16_MPORT_data = rf[rf_io_dbg_monitor_reg_16_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_17_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_17_MPORT_addr = 5'h11;
  assign rf_io_dbg_monitor_reg_17_MPORT_data = rf[rf_io_dbg_monitor_reg_17_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_18_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_18_MPORT_addr = 5'h12;
  assign rf_io_dbg_monitor_reg_18_MPORT_data = rf[rf_io_dbg_monitor_reg_18_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_19_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_19_MPORT_addr = 5'h13;
  assign rf_io_dbg_monitor_reg_19_MPORT_data = rf[rf_io_dbg_monitor_reg_19_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_20_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_20_MPORT_addr = 5'h14;
  assign rf_io_dbg_monitor_reg_20_MPORT_data = rf[rf_io_dbg_monitor_reg_20_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_21_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_21_MPORT_addr = 5'h15;
  assign rf_io_dbg_monitor_reg_21_MPORT_data = rf[rf_io_dbg_monitor_reg_21_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_22_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_22_MPORT_addr = 5'h16;
  assign rf_io_dbg_monitor_reg_22_MPORT_data = rf[rf_io_dbg_monitor_reg_22_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_23_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_23_MPORT_addr = 5'h17;
  assign rf_io_dbg_monitor_reg_23_MPORT_data = rf[rf_io_dbg_monitor_reg_23_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_24_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_24_MPORT_addr = 5'h18;
  assign rf_io_dbg_monitor_reg_24_MPORT_data = rf[rf_io_dbg_monitor_reg_24_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_25_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_25_MPORT_addr = 5'h19;
  assign rf_io_dbg_monitor_reg_25_MPORT_data = rf[rf_io_dbg_monitor_reg_25_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_26_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_26_MPORT_addr = 5'h1a;
  assign rf_io_dbg_monitor_reg_26_MPORT_data = rf[rf_io_dbg_monitor_reg_26_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_27_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_27_MPORT_addr = 5'h1b;
  assign rf_io_dbg_monitor_reg_27_MPORT_data = rf[rf_io_dbg_monitor_reg_27_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_28_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_28_MPORT_addr = 5'h1c;
  assign rf_io_dbg_monitor_reg_28_MPORT_data = rf[rf_io_dbg_monitor_reg_28_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_29_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_29_MPORT_addr = 5'h1d;
  assign rf_io_dbg_monitor_reg_29_MPORT_data = rf[rf_io_dbg_monitor_reg_29_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_30_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_30_MPORT_addr = 5'h1e;
  assign rf_io_dbg_monitor_reg_30_MPORT_data = rf[rf_io_dbg_monitor_reg_30_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_io_dbg_monitor_reg_31_MPORT_en = 1'h1;
  assign rf_io_dbg_monitor_reg_31_MPORT_addr = 5'h1f;
  assign rf_io_dbg_monitor_reg_31_MPORT_data = rf[rf_io_dbg_monitor_reg_31_MPORT_addr]; // @[Register.scala 8:15]
  assign rf_MPORT_data = wb_ctrl_jalr ? wb_npc : _rf_wdata_T_4;
  assign rf_MPORT_addr = wb_reg_waddr;
  assign rf_MPORT_mask = 1'h1;
  assign rf_MPORT_en = wb_ctrl_wxd & _T_7;
  assign io_iData_addr = pc; // @[RISCV.scala 137:17]
  assign io_dData_addr = mem_alu_out; // @[RISCV.scala 331:17]
  assign io_dData_writeData = mem_rs_1; // @[RISCV.scala 337:22]
  assign io_dData_writeEnable = mem_ctrl_mem_cmd == 5'h1; // @[RISCV.scala 333:44]
  assign alu_io_fn = ex_ctrl_alu_fn; // @[RISCV.scala 290:13]
  assign alu_io_in1 = 2'h2 == ex_ctrl_sel_alu1 ? ex_pc : _ex_op1_T_1; // @[Mux.scala 81:58]
  assign alu_io_in2 = 2'h1 == ex_ctrl_sel_alu2 ? 32'h4 : _ex_op2_T_4; // @[Mux.scala 81:58]
  assign rf_clock = ~clock;
  always @(posedge rf_clock) begin
    if (rf_MPORT_en & rf_MPORT_mask) begin
      rf[rf_MPORT_addr] <= rf_MPORT_data; // @[Register.scala 8:15]
    end
  end
  always @(posedge clock) begin
    if (reset) begin // @[RISCV.scala 58:22]
      id_pc <= 32'h80000000; // @[RISCV.scala 58:22]
    end else if (~load_stall & ~jump_flush) begin // @[RISCV.scala 152:36]
      id_pc <= pc; // @[RISCV.scala 153:11]
    end else if (jump_flush) begin // @[RISCV.scala 156:26]
      id_pc <= 32'h80000000; // @[RISCV.scala 157:11]
    end
    if (reset) begin // @[RISCV.scala 59:23]
      id_npc <= 32'h80000004; // @[RISCV.scala 59:23]
    end else if (~load_stall & ~jump_flush) begin // @[RISCV.scala 152:36]
      id_npc <= npc; // @[RISCV.scala 154:12]
    end else if (jump_flush) begin // @[RISCV.scala 156:26]
      id_npc <= 32'h80000004; // @[RISCV.scala 158:12]
    end
    if (reset) begin // @[RISCV.scala 60:24]
      id_inst <= 32'h13; // @[RISCV.scala 60:24]
    end else if (~load_stall & ~jump_flush) begin // @[RISCV.scala 152:36]
      id_inst <= io_iData_inst; // @[RISCV.scala 155:13]
    end else if (jump_flush) begin // @[RISCV.scala 156:26]
      id_inst <= 32'h13; // @[RISCV.scala 159:13]
    end
    if (reset) begin // @[RISCV.scala 70:22]
      ex_pc <= 32'h80000000; // @[RISCV.scala 70:22]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_pc <= id_pc; // @[RISCV.scala 213:11]
    end else begin
      ex_pc <= 32'h80000000; // @[RISCV.scala 221:11]
    end
    if (reset) begin // @[RISCV.scala 71:23]
      ex_npc <= 32'h80000004; // @[RISCV.scala 71:23]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_npc <= id_npc; // @[RISCV.scala 214:12]
    end else begin
      ex_npc <= 32'h80000004; // @[RISCV.scala 222:12]
    end
    if (reset) begin // @[RISCV.scala 72:24]
      ex_inst <= 32'h13; // @[RISCV.scala 72:24]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_inst <= id_inst; // @[RISCV.scala 215:13]
    end else begin
      ex_inst <= 32'h13; // @[RISCV.scala 224:13]
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_branch <= 1'h0; // @[RISCV.scala 73:24]
    end else begin
      ex_ctrl_branch <= _GEN_19;
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_jal <= 1'h0; // @[RISCV.scala 73:24]
    end else begin
      ex_ctrl_jal <= _GEN_18;
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_jalr <= 1'h0; // @[RISCV.scala 73:24]
    end else begin
      ex_ctrl_jalr <= _GEN_17;
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_sel_alu1 <= 2'h1; // @[RISCV.scala 73:24]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      if (id_ctrl_decoder_0) begin // @[Mux.scala 101:16]
        ex_ctrl_sel_alu1 <= 2'h1;
      end else if (_id_ctrl_decoder_ctrl_signals_T_3) begin // @[Mux.scala 101:16]
        ex_ctrl_sel_alu1 <= 2'h1;
      end else begin
        ex_ctrl_sel_alu1 <= _id_ctrl_decoder_ctrl_signals_T_90;
      end
    end else begin
      ex_ctrl_sel_alu1 <= 2'h1; // @[RISCV.scala 223:13]
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_sel_alu2 <= 2'h3; // @[RISCV.scala 73:24]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      if (id_ctrl_decoder_0) begin // @[Mux.scala 101:16]
        ex_ctrl_sel_alu2 <= 2'h2;
      end else if (_id_ctrl_decoder_ctrl_signals_T_3) begin // @[Mux.scala 101:16]
        ex_ctrl_sel_alu2 <= 2'h3;
      end else begin
        ex_ctrl_sel_alu2 <= _id_ctrl_decoder_ctrl_signals_T_113;
      end
    end else begin
      ex_ctrl_sel_alu2 <= 2'h3; // @[RISCV.scala 223:13]
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_sel_imm <= 3'h4; // @[RISCV.scala 73:24]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      if (id_ctrl_decoder_0) begin // @[Mux.scala 101:16]
        ex_ctrl_sel_imm <= 3'h1;
      end else if (_id_ctrl_decoder_ctrl_signals_T_3) begin // @[Mux.scala 101:16]
        ex_ctrl_sel_imm <= 3'h4;
      end else begin
        ex_ctrl_sel_imm <= _id_ctrl_decoder_ctrl_signals_T_136;
      end
    end else begin
      ex_ctrl_sel_imm <= 3'h4; // @[RISCV.scala 223:13]
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_alu_fn <= 4'h0; // @[RISCV.scala 73:24]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_ctrl_alu_fn <= id_ctrl_alu_fn; // @[RISCV.scala 216:13]
    end else begin
      ex_ctrl_alu_fn <= 4'h0; // @[RISCV.scala 223:13]
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_mem <= 1'h0; // @[RISCV.scala 73:24]
    end else begin
      ex_ctrl_mem <= _GEN_12;
    end
    if (reset) begin // @[RISCV.scala 73:24]
      ex_ctrl_mem_cmd <= 5'h0; // @[RISCV.scala 73:24]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_ctrl_mem_cmd <= id_ctrl_mem_cmd; // @[RISCV.scala 216:13]
    end else begin
      ex_ctrl_mem_cmd <= 5'h0; // @[RISCV.scala 223:13]
    end
    ex_ctrl_wxd <= reset | _GEN_9; // @[RISCV.scala 73:{24,24}]
    if (reset) begin // @[RISCV.scala 74:29]
      ex_reg_raddr_0 <= 5'h0; // @[RISCV.scala 74:29]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_reg_raddr_0 <= id_inst_arange_rs1; // @[RISCV.scala 217:18]
    end else begin
      ex_reg_raddr_0 <= 5'h0; // @[RISCV.scala 225:18]
    end
    if (reset) begin // @[RISCV.scala 74:29]
      ex_reg_raddr_1 <= 5'h0; // @[RISCV.scala 74:29]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_reg_raddr_1 <= id_inst_arange_rs2; // @[RISCV.scala 217:18]
    end else begin
      ex_reg_raddr_1 <= 5'h0; // @[RISCV.scala 225:18]
    end
    if (reset) begin // @[RISCV.scala 75:29]
      ex_reg_waddr <= 5'h0; // @[RISCV.scala 75:29]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      ex_reg_waddr <= id_inst_arange_rd; // @[RISCV.scala 218:18]
    end else begin
      ex_reg_waddr <= 5'h0; // @[RISCV.scala 226:18]
    end
    if (reset) begin // @[RISCV.scala 76:22]
      ex_rs_0 <= 32'h0; // @[RISCV.scala 76:22]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      if (id_inst_arange_rs1 == 5'h0) begin // @[Register.scala 12:8]
        ex_rs_0 <= 32'h0;
      end else begin
        ex_rs_0 <= rf_id_rs_MPORT_data;
      end
    end else begin
      ex_rs_0 <= 32'h0; // @[RISCV.scala 227:11]
    end
    if (reset) begin // @[RISCV.scala 76:22]
      ex_rs_1 <= 32'h0; // @[RISCV.scala 76:22]
    end else if (_T_2) begin // @[RISCV.scala 212:36]
      if (id_inst_arange_rs2 == 5'h0) begin // @[Register.scala 12:8]
        ex_rs_1 <= 32'h0;
      end else begin
        ex_rs_1 <= rf_id_rs_MPORT_1_data;
      end
    end else begin
      ex_rs_1 <= 32'h0; // @[RISCV.scala 227:11]
    end
    if (reset) begin // @[RISCV.scala 87:23]
      mem_pc <= 32'h80000000; // @[RISCV.scala 87:23]
    end else if (_T_1) begin // @[RISCV.scala 308:21]
      mem_pc <= ex_pc; // @[RISCV.scala 309:12]
    end else begin
      mem_pc <= 32'h80000000; // @[RISCV.scala 318:12]
    end
    if (reset) begin // @[RISCV.scala 88:24]
      mem_npc <= 32'h80000004; // @[RISCV.scala 88:24]
    end else if (_T_1) begin // @[RISCV.scala 308:21]
      mem_npc <= ex_npc; // @[RISCV.scala 310:13]
    end else begin
      mem_npc <= 32'h80000004; // @[RISCV.scala 319:13]
    end
    if (reset) begin // @[RISCV.scala 89:25]
      mem_ctrl_branch <= 1'h0; // @[RISCV.scala 89:25]
    end else begin
      mem_ctrl_branch <= _GEN_37;
    end
    if (reset) begin // @[RISCV.scala 89:25]
      mem_ctrl_jal <= 1'h0; // @[RISCV.scala 89:25]
    end else begin
      mem_ctrl_jal <= _GEN_36;
    end
    if (reset) begin // @[RISCV.scala 89:25]
      mem_ctrl_jalr <= 1'h0; // @[RISCV.scala 89:25]
    end else begin
      mem_ctrl_jalr <= _GEN_35;
    end
    if (reset) begin // @[RISCV.scala 89:25]
      mem_ctrl_mem <= 1'h0; // @[RISCV.scala 89:25]
    end else begin
      mem_ctrl_mem <= _GEN_30;
    end
    if (reset) begin // @[RISCV.scala 89:25]
      mem_ctrl_mem_cmd <= 5'h0; // @[RISCV.scala 89:25]
    end else if (_T_1) begin // @[RISCV.scala 308:21]
      mem_ctrl_mem_cmd <= ex_ctrl_mem_cmd; // @[RISCV.scala 311:14]
    end else begin
      mem_ctrl_mem_cmd <= 5'h0; // @[RISCV.scala 320:14]
    end
    mem_ctrl_wxd <= reset | _GEN_27; // @[RISCV.scala 89:{25,25}]
    if (reset) begin // @[RISCV.scala 90:30]
      mem_reg_waddr <= 5'h0; // @[RISCV.scala 90:30]
    end else if (_T_1) begin // @[RISCV.scala 308:21]
      mem_reg_waddr <= ex_reg_waddr; // @[RISCV.scala 313:19]
    end else begin
      mem_reg_waddr <= 5'h0; // @[RISCV.scala 322:19]
    end
    if (reset) begin // @[RISCV.scala 91:23]
      mem_rs_1 <= 32'h0; // @[RISCV.scala 91:23]
    end else if (_T_1) begin // @[RISCV.scala 308:21]
      if (_ex_rs_bypassed_T_21) begin // @[Mux.scala 101:16]
        mem_rs_1 <= mem_alu_out;
      end else if (_ex_rs_bypassed_T_30) begin // @[Mux.scala 101:16]
        mem_rs_1 <= io_dData_readData;
      end else begin
        mem_rs_1 <= ex_rs_1;
      end
    end else begin
      mem_rs_1 <= 32'h0; // @[RISCV.scala 321:12]
    end
    if (reset) begin // @[RISCV.scala 92:24]
      mem_imm <= 32'sh0; // @[RISCV.scala 92:24]
    end else if (_T_1) begin // @[RISCV.scala 308:21]
      mem_imm <= ex_imm; // @[RISCV.scala 314:13]
    end else begin
      mem_imm <= 32'sh0; // @[RISCV.scala 323:13]
    end
    if (reset) begin // @[RISCV.scala 93:28]
      mem_alu_out <= 32'h0; // @[RISCV.scala 93:28]
    end else if (_T_1) begin // @[RISCV.scala 308:21]
      mem_alu_out <= alu_io_alu_out; // @[RISCV.scala 315:17]
    end else begin
      mem_alu_out <= 32'h0; // @[RISCV.scala 324:17]
    end
    if (reset) begin // @[RISCV.scala 94:32]
      mem_alu_cmp_out <= 1'h0; // @[RISCV.scala 94:32]
    end else begin
      mem_alu_cmp_out <= _GEN_43;
    end
    if (reset) begin // @[RISCV.scala 102:23]
      wb_npc <= 32'h80000004; // @[RISCV.scala 102:23]
    end else begin
      wb_npc <= mem_npc; // @[RISCV.scala 349:10]
    end
    if (reset) begin // @[RISCV.scala 103:24]
      wb_ctrl_jalr <= 1'h0; // @[RISCV.scala 103:24]
    end else begin
      wb_ctrl_jalr <= mem_ctrl_jalr; // @[RISCV.scala 350:11]
    end
    if (reset) begin // @[RISCV.scala 103:24]
      wb_ctrl_mem <= 1'h0; // @[RISCV.scala 103:24]
    end else begin
      wb_ctrl_mem <= mem_ctrl_mem; // @[RISCV.scala 350:11]
    end
    wb_ctrl_wxd <= reset | mem_ctrl_wxd; // @[RISCV.scala 103:{24,24} 350:11]
    if (reset) begin // @[RISCV.scala 105:29]
      wb_reg_waddr <= 5'h0; // @[RISCV.scala 105:29]
    end else begin
      wb_reg_waddr <= mem_reg_waddr; // @[RISCV.scala 351:16]
    end
    if (reset) begin // @[RISCV.scala 106:27]
      wb_alu_out <= 32'h0; // @[RISCV.scala 106:27]
    end else begin
      wb_alu_out <= mem_alu_out; // @[RISCV.scala 352:14]
    end
    if (reset) begin // @[RISCV.scala 107:34]
      wb_dData_readData <= 32'h0; // @[RISCV.scala 107:34]
    end else begin
      wb_dData_readData <= io_dData_readData; // @[RISCV.scala 353:21]
    end
    if (reset) begin // @[RISCV.scala 127:19]
      pc <= 32'h80000000; // @[RISCV.scala 127:19]
    end else if (_T) begin // @[RISCV.scala 380:21]
      if (_jump_flush_T_5) begin // @[Mux.scala 101:16]
        pc <= _pc_T_8;
      end else if (mem_ctrl_jalr) begin // @[Mux.scala 101:16]
        pc <= mem_alu_out;
      end else begin
        pc <= npc;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    rf[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  id_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  id_npc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  id_inst = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  ex_pc = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  ex_npc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  ex_inst = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ex_ctrl_branch = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  ex_ctrl_jal = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  ex_ctrl_jalr = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ex_ctrl_sel_alu1 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  ex_ctrl_sel_alu2 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  ex_ctrl_sel_imm = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  ex_ctrl_alu_fn = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  ex_ctrl_mem = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ex_ctrl_mem_cmd = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  ex_ctrl_wxd = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ex_reg_raddr_0 = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  ex_reg_raddr_1 = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  ex_reg_waddr = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  ex_rs_0 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  ex_rs_1 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mem_pc = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mem_npc = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  mem_ctrl_branch = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  mem_ctrl_jal = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  mem_ctrl_jalr = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  mem_ctrl_mem = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  mem_ctrl_mem_cmd = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  mem_ctrl_wxd = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  mem_reg_waddr = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  mem_rs_1 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  mem_imm = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  mem_alu_out = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  mem_alu_cmp_out = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  wb_npc = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  wb_ctrl_jalr = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  wb_ctrl_mem = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  wb_ctrl_wxd = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  wb_reg_waddr = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  wb_alu_out = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  wb_dData_readData = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  pc = _RAND_42[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IData(
  input  [31:0] io_addr,
  output [31:0] io_inst
);
  wire [31:0] _GEN_1 = 8'h1 == io_addr[9:2] ? 32'h2c40413 : 32'h417; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_2 = 8'h2 == io_addr[9:2] ? 32'h40503 : _GEN_1; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_3 = 8'h3 == io_addr[9:2] ? 32'h140413 : _GEN_2; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_4 = 8'h4 == io_addr[9:2] ? 32'h50c63 : _GEN_3; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_5 = 8'h5 == io_addr[9:2] ? 32'h8000ef : _GEN_4; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_6 = 8'h6 == io_addr[9:2] ? 32'hff1ff06f : _GEN_5; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_7 = 8'h7 == io_addr[9:2] ? 32'h100002b7 : _GEN_6; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_8 = 8'h8 == io_addr[9:2] ? 32'ha28023 : _GEN_7; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_9 = 8'h9 == io_addr[9:2] ? 32'h8067 : _GEN_8; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_10 = 8'ha == io_addr[9:2] ? 32'h6f : _GEN_9; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_11 = 8'hb == io_addr[9:2] ? 32'h0 : _GEN_10; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_12 = 8'hc == io_addr[9:2] ? 32'h0 : _GEN_11; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_13 = 8'hd == io_addr[9:2] ? 32'h0 : _GEN_12; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_14 = 8'he == io_addr[9:2] ? 32'h0 : _GEN_13; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_15 = 8'hf == io_addr[9:2] ? 32'h0 : _GEN_14; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_16 = 8'h10 == io_addr[9:2] ? 32'h0 : _GEN_15; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_17 = 8'h11 == io_addr[9:2] ? 32'h0 : _GEN_16; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_18 = 8'h12 == io_addr[9:2] ? 32'h0 : _GEN_17; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_19 = 8'h13 == io_addr[9:2] ? 32'h0 : _GEN_18; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_20 = 8'h14 == io_addr[9:2] ? 32'h0 : _GEN_19; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_21 = 8'h15 == io_addr[9:2] ? 32'h0 : _GEN_20; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_22 = 8'h16 == io_addr[9:2] ? 32'h0 : _GEN_21; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_23 = 8'h17 == io_addr[9:2] ? 32'h0 : _GEN_22; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_24 = 8'h18 == io_addr[9:2] ? 32'h0 : _GEN_23; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_25 = 8'h19 == io_addr[9:2] ? 32'h0 : _GEN_24; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_26 = 8'h1a == io_addr[9:2] ? 32'h0 : _GEN_25; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_27 = 8'h1b == io_addr[9:2] ? 32'h0 : _GEN_26; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_28 = 8'h1c == io_addr[9:2] ? 32'h0 : _GEN_27; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_29 = 8'h1d == io_addr[9:2] ? 32'h0 : _GEN_28; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_30 = 8'h1e == io_addr[9:2] ? 32'h0 : _GEN_29; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_31 = 8'h1f == io_addr[9:2] ? 32'h0 : _GEN_30; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_32 = 8'h20 == io_addr[9:2] ? 32'h0 : _GEN_31; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_33 = 8'h21 == io_addr[9:2] ? 32'h0 : _GEN_32; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_34 = 8'h22 == io_addr[9:2] ? 32'h0 : _GEN_33; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_35 = 8'h23 == io_addr[9:2] ? 32'h0 : _GEN_34; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_36 = 8'h24 == io_addr[9:2] ? 32'h0 : _GEN_35; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_37 = 8'h25 == io_addr[9:2] ? 32'h0 : _GEN_36; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_38 = 8'h26 == io_addr[9:2] ? 32'h0 : _GEN_37; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_39 = 8'h27 == io_addr[9:2] ? 32'h0 : _GEN_38; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_40 = 8'h28 == io_addr[9:2] ? 32'h0 : _GEN_39; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_41 = 8'h29 == io_addr[9:2] ? 32'h0 : _GEN_40; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_42 = 8'h2a == io_addr[9:2] ? 32'h0 : _GEN_41; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_43 = 8'h2b == io_addr[9:2] ? 32'h0 : _GEN_42; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_44 = 8'h2c == io_addr[9:2] ? 32'h0 : _GEN_43; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_45 = 8'h2d == io_addr[9:2] ? 32'h0 : _GEN_44; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_46 = 8'h2e == io_addr[9:2] ? 32'h0 : _GEN_45; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_47 = 8'h2f == io_addr[9:2] ? 32'h0 : _GEN_46; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_48 = 8'h30 == io_addr[9:2] ? 32'h0 : _GEN_47; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_49 = 8'h31 == io_addr[9:2] ? 32'h0 : _GEN_48; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_50 = 8'h32 == io_addr[9:2] ? 32'h0 : _GEN_49; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_51 = 8'h33 == io_addr[9:2] ? 32'h0 : _GEN_50; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_52 = 8'h34 == io_addr[9:2] ? 32'h0 : _GEN_51; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_53 = 8'h35 == io_addr[9:2] ? 32'h0 : _GEN_52; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_54 = 8'h36 == io_addr[9:2] ? 32'h0 : _GEN_53; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_55 = 8'h37 == io_addr[9:2] ? 32'h0 : _GEN_54; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_56 = 8'h38 == io_addr[9:2] ? 32'h0 : _GEN_55; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_57 = 8'h39 == io_addr[9:2] ? 32'h0 : _GEN_56; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_58 = 8'h3a == io_addr[9:2] ? 32'h0 : _GEN_57; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_59 = 8'h3b == io_addr[9:2] ? 32'h0 : _GEN_58; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_60 = 8'h3c == io_addr[9:2] ? 32'h0 : _GEN_59; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_61 = 8'h3d == io_addr[9:2] ? 32'h0 : _GEN_60; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_62 = 8'h3e == io_addr[9:2] ? 32'h0 : _GEN_61; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_63 = 8'h3f == io_addr[9:2] ? 32'h0 : _GEN_62; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_64 = 8'h40 == io_addr[9:2] ? 32'h0 : _GEN_63; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_65 = 8'h41 == io_addr[9:2] ? 32'h0 : _GEN_64; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_66 = 8'h42 == io_addr[9:2] ? 32'h0 : _GEN_65; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_67 = 8'h43 == io_addr[9:2] ? 32'h0 : _GEN_66; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_68 = 8'h44 == io_addr[9:2] ? 32'h0 : _GEN_67; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_69 = 8'h45 == io_addr[9:2] ? 32'h0 : _GEN_68; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_70 = 8'h46 == io_addr[9:2] ? 32'h0 : _GEN_69; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_71 = 8'h47 == io_addr[9:2] ? 32'h0 : _GEN_70; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_72 = 8'h48 == io_addr[9:2] ? 32'h0 : _GEN_71; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_73 = 8'h49 == io_addr[9:2] ? 32'h0 : _GEN_72; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_74 = 8'h4a == io_addr[9:2] ? 32'h0 : _GEN_73; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_75 = 8'h4b == io_addr[9:2] ? 32'h0 : _GEN_74; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_76 = 8'h4c == io_addr[9:2] ? 32'h0 : _GEN_75; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_77 = 8'h4d == io_addr[9:2] ? 32'h0 : _GEN_76; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_78 = 8'h4e == io_addr[9:2] ? 32'h0 : _GEN_77; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_79 = 8'h4f == io_addr[9:2] ? 32'h0 : _GEN_78; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_80 = 8'h50 == io_addr[9:2] ? 32'h0 : _GEN_79; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_81 = 8'h51 == io_addr[9:2] ? 32'h0 : _GEN_80; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_82 = 8'h52 == io_addr[9:2] ? 32'h0 : _GEN_81; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_83 = 8'h53 == io_addr[9:2] ? 32'h0 : _GEN_82; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_84 = 8'h54 == io_addr[9:2] ? 32'h0 : _GEN_83; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_85 = 8'h55 == io_addr[9:2] ? 32'h0 : _GEN_84; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_86 = 8'h56 == io_addr[9:2] ? 32'h0 : _GEN_85; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_87 = 8'h57 == io_addr[9:2] ? 32'h0 : _GEN_86; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_88 = 8'h58 == io_addr[9:2] ? 32'h0 : _GEN_87; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_89 = 8'h59 == io_addr[9:2] ? 32'h0 : _GEN_88; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_90 = 8'h5a == io_addr[9:2] ? 32'h0 : _GEN_89; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_91 = 8'h5b == io_addr[9:2] ? 32'h0 : _GEN_90; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_92 = 8'h5c == io_addr[9:2] ? 32'h0 : _GEN_91; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_93 = 8'h5d == io_addr[9:2] ? 32'h0 : _GEN_92; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_94 = 8'h5e == io_addr[9:2] ? 32'h0 : _GEN_93; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_95 = 8'h5f == io_addr[9:2] ? 32'h0 : _GEN_94; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_96 = 8'h60 == io_addr[9:2] ? 32'h0 : _GEN_95; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_97 = 8'h61 == io_addr[9:2] ? 32'h0 : _GEN_96; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_98 = 8'h62 == io_addr[9:2] ? 32'h0 : _GEN_97; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_99 = 8'h63 == io_addr[9:2] ? 32'h0 : _GEN_98; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_100 = 8'h64 == io_addr[9:2] ? 32'h0 : _GEN_99; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_101 = 8'h65 == io_addr[9:2] ? 32'h0 : _GEN_100; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_102 = 8'h66 == io_addr[9:2] ? 32'h0 : _GEN_101; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_103 = 8'h67 == io_addr[9:2] ? 32'h0 : _GEN_102; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_104 = 8'h68 == io_addr[9:2] ? 32'h0 : _GEN_103; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_105 = 8'h69 == io_addr[9:2] ? 32'h0 : _GEN_104; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_106 = 8'h6a == io_addr[9:2] ? 32'h0 : _GEN_105; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_107 = 8'h6b == io_addr[9:2] ? 32'h0 : _GEN_106; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_108 = 8'h6c == io_addr[9:2] ? 32'h0 : _GEN_107; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_109 = 8'h6d == io_addr[9:2] ? 32'h0 : _GEN_108; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_110 = 8'h6e == io_addr[9:2] ? 32'h0 : _GEN_109; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_111 = 8'h6f == io_addr[9:2] ? 32'h0 : _GEN_110; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_112 = 8'h70 == io_addr[9:2] ? 32'h0 : _GEN_111; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_113 = 8'h71 == io_addr[9:2] ? 32'h0 : _GEN_112; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_114 = 8'h72 == io_addr[9:2] ? 32'h0 : _GEN_113; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_115 = 8'h73 == io_addr[9:2] ? 32'h0 : _GEN_114; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_116 = 8'h74 == io_addr[9:2] ? 32'h0 : _GEN_115; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_117 = 8'h75 == io_addr[9:2] ? 32'h0 : _GEN_116; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_118 = 8'h76 == io_addr[9:2] ? 32'h0 : _GEN_117; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_119 = 8'h77 == io_addr[9:2] ? 32'h0 : _GEN_118; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_120 = 8'h78 == io_addr[9:2] ? 32'h0 : _GEN_119; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_121 = 8'h79 == io_addr[9:2] ? 32'h0 : _GEN_120; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_122 = 8'h7a == io_addr[9:2] ? 32'h0 : _GEN_121; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_123 = 8'h7b == io_addr[9:2] ? 32'h0 : _GEN_122; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_124 = 8'h7c == io_addr[9:2] ? 32'h0 : _GEN_123; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_125 = 8'h7d == io_addr[9:2] ? 32'h0 : _GEN_124; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_126 = 8'h7e == io_addr[9:2] ? 32'h0 : _GEN_125; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_127 = 8'h7f == io_addr[9:2] ? 32'h0 : _GEN_126; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_128 = 8'h80 == io_addr[9:2] ? 32'h0 : _GEN_127; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_129 = 8'h81 == io_addr[9:2] ? 32'h0 : _GEN_128; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_130 = 8'h82 == io_addr[9:2] ? 32'h0 : _GEN_129; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_131 = 8'h83 == io_addr[9:2] ? 32'h0 : _GEN_130; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_132 = 8'h84 == io_addr[9:2] ? 32'h0 : _GEN_131; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_133 = 8'h85 == io_addr[9:2] ? 32'h0 : _GEN_132; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_134 = 8'h86 == io_addr[9:2] ? 32'h0 : _GEN_133; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_135 = 8'h87 == io_addr[9:2] ? 32'h0 : _GEN_134; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_136 = 8'h88 == io_addr[9:2] ? 32'h0 : _GEN_135; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_137 = 8'h89 == io_addr[9:2] ? 32'h0 : _GEN_136; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_138 = 8'h8a == io_addr[9:2] ? 32'h0 : _GEN_137; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_139 = 8'h8b == io_addr[9:2] ? 32'h0 : _GEN_138; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_140 = 8'h8c == io_addr[9:2] ? 32'h0 : _GEN_139; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_141 = 8'h8d == io_addr[9:2] ? 32'h0 : _GEN_140; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_142 = 8'h8e == io_addr[9:2] ? 32'h0 : _GEN_141; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_143 = 8'h8f == io_addr[9:2] ? 32'h0 : _GEN_142; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_144 = 8'h90 == io_addr[9:2] ? 32'h0 : _GEN_143; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_145 = 8'h91 == io_addr[9:2] ? 32'h0 : _GEN_144; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_146 = 8'h92 == io_addr[9:2] ? 32'h0 : _GEN_145; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_147 = 8'h93 == io_addr[9:2] ? 32'h0 : _GEN_146; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_148 = 8'h94 == io_addr[9:2] ? 32'h0 : _GEN_147; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_149 = 8'h95 == io_addr[9:2] ? 32'h0 : _GEN_148; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_150 = 8'h96 == io_addr[9:2] ? 32'h0 : _GEN_149; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_151 = 8'h97 == io_addr[9:2] ? 32'h0 : _GEN_150; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_152 = 8'h98 == io_addr[9:2] ? 32'h0 : _GEN_151; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_153 = 8'h99 == io_addr[9:2] ? 32'h0 : _GEN_152; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_154 = 8'h9a == io_addr[9:2] ? 32'h0 : _GEN_153; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_155 = 8'h9b == io_addr[9:2] ? 32'h0 : _GEN_154; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_156 = 8'h9c == io_addr[9:2] ? 32'h0 : _GEN_155; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_157 = 8'h9d == io_addr[9:2] ? 32'h0 : _GEN_156; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_158 = 8'h9e == io_addr[9:2] ? 32'h0 : _GEN_157; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_159 = 8'h9f == io_addr[9:2] ? 32'h0 : _GEN_158; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_160 = 8'ha0 == io_addr[9:2] ? 32'h0 : _GEN_159; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_161 = 8'ha1 == io_addr[9:2] ? 32'h0 : _GEN_160; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_162 = 8'ha2 == io_addr[9:2] ? 32'h0 : _GEN_161; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_163 = 8'ha3 == io_addr[9:2] ? 32'h0 : _GEN_162; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_164 = 8'ha4 == io_addr[9:2] ? 32'h0 : _GEN_163; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_165 = 8'ha5 == io_addr[9:2] ? 32'h0 : _GEN_164; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_166 = 8'ha6 == io_addr[9:2] ? 32'h0 : _GEN_165; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_167 = 8'ha7 == io_addr[9:2] ? 32'h0 : _GEN_166; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_168 = 8'ha8 == io_addr[9:2] ? 32'h0 : _GEN_167; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_169 = 8'ha9 == io_addr[9:2] ? 32'h0 : _GEN_168; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_170 = 8'haa == io_addr[9:2] ? 32'h0 : _GEN_169; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_171 = 8'hab == io_addr[9:2] ? 32'h0 : _GEN_170; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_172 = 8'hac == io_addr[9:2] ? 32'h0 : _GEN_171; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_173 = 8'had == io_addr[9:2] ? 32'h0 : _GEN_172; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_174 = 8'hae == io_addr[9:2] ? 32'h0 : _GEN_173; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_175 = 8'haf == io_addr[9:2] ? 32'h0 : _GEN_174; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_176 = 8'hb0 == io_addr[9:2] ? 32'h0 : _GEN_175; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_177 = 8'hb1 == io_addr[9:2] ? 32'h0 : _GEN_176; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_178 = 8'hb2 == io_addr[9:2] ? 32'h0 : _GEN_177; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_179 = 8'hb3 == io_addr[9:2] ? 32'h0 : _GEN_178; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_180 = 8'hb4 == io_addr[9:2] ? 32'h0 : _GEN_179; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_181 = 8'hb5 == io_addr[9:2] ? 32'h0 : _GEN_180; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_182 = 8'hb6 == io_addr[9:2] ? 32'h0 : _GEN_181; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_183 = 8'hb7 == io_addr[9:2] ? 32'h0 : _GEN_182; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_184 = 8'hb8 == io_addr[9:2] ? 32'h0 : _GEN_183; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_185 = 8'hb9 == io_addr[9:2] ? 32'h0 : _GEN_184; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_186 = 8'hba == io_addr[9:2] ? 32'h0 : _GEN_185; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_187 = 8'hbb == io_addr[9:2] ? 32'h0 : _GEN_186; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_188 = 8'hbc == io_addr[9:2] ? 32'h0 : _GEN_187; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_189 = 8'hbd == io_addr[9:2] ? 32'h0 : _GEN_188; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_190 = 8'hbe == io_addr[9:2] ? 32'h0 : _GEN_189; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_191 = 8'hbf == io_addr[9:2] ? 32'h0 : _GEN_190; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_192 = 8'hc0 == io_addr[9:2] ? 32'h0 : _GEN_191; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_193 = 8'hc1 == io_addr[9:2] ? 32'h0 : _GEN_192; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_194 = 8'hc2 == io_addr[9:2] ? 32'h0 : _GEN_193; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_195 = 8'hc3 == io_addr[9:2] ? 32'h0 : _GEN_194; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_196 = 8'hc4 == io_addr[9:2] ? 32'h0 : _GEN_195; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_197 = 8'hc5 == io_addr[9:2] ? 32'h0 : _GEN_196; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_198 = 8'hc6 == io_addr[9:2] ? 32'h0 : _GEN_197; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_199 = 8'hc7 == io_addr[9:2] ? 32'h0 : _GEN_198; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_200 = 8'hc8 == io_addr[9:2] ? 32'h0 : _GEN_199; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_201 = 8'hc9 == io_addr[9:2] ? 32'h0 : _GEN_200; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_202 = 8'hca == io_addr[9:2] ? 32'h0 : _GEN_201; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_203 = 8'hcb == io_addr[9:2] ? 32'h0 : _GEN_202; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_204 = 8'hcc == io_addr[9:2] ? 32'h0 : _GEN_203; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_205 = 8'hcd == io_addr[9:2] ? 32'h0 : _GEN_204; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_206 = 8'hce == io_addr[9:2] ? 32'h0 : _GEN_205; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_207 = 8'hcf == io_addr[9:2] ? 32'h0 : _GEN_206; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_208 = 8'hd0 == io_addr[9:2] ? 32'h0 : _GEN_207; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_209 = 8'hd1 == io_addr[9:2] ? 32'h0 : _GEN_208; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_210 = 8'hd2 == io_addr[9:2] ? 32'h0 : _GEN_209; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_211 = 8'hd3 == io_addr[9:2] ? 32'h0 : _GEN_210; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_212 = 8'hd4 == io_addr[9:2] ? 32'h0 : _GEN_211; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_213 = 8'hd5 == io_addr[9:2] ? 32'h0 : _GEN_212; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_214 = 8'hd6 == io_addr[9:2] ? 32'h0 : _GEN_213; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_215 = 8'hd7 == io_addr[9:2] ? 32'h0 : _GEN_214; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_216 = 8'hd8 == io_addr[9:2] ? 32'h0 : _GEN_215; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_217 = 8'hd9 == io_addr[9:2] ? 32'h0 : _GEN_216; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_218 = 8'hda == io_addr[9:2] ? 32'h0 : _GEN_217; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_219 = 8'hdb == io_addr[9:2] ? 32'h0 : _GEN_218; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_220 = 8'hdc == io_addr[9:2] ? 32'h0 : _GEN_219; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_221 = 8'hdd == io_addr[9:2] ? 32'h0 : _GEN_220; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_222 = 8'hde == io_addr[9:2] ? 32'h0 : _GEN_221; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_223 = 8'hdf == io_addr[9:2] ? 32'h0 : _GEN_222; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_224 = 8'he0 == io_addr[9:2] ? 32'h0 : _GEN_223; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_225 = 8'he1 == io_addr[9:2] ? 32'h0 : _GEN_224; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_226 = 8'he2 == io_addr[9:2] ? 32'h0 : _GEN_225; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_227 = 8'he3 == io_addr[9:2] ? 32'h0 : _GEN_226; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_228 = 8'he4 == io_addr[9:2] ? 32'h0 : _GEN_227; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_229 = 8'he5 == io_addr[9:2] ? 32'h0 : _GEN_228; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_230 = 8'he6 == io_addr[9:2] ? 32'h0 : _GEN_229; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_231 = 8'he7 == io_addr[9:2] ? 32'h0 : _GEN_230; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_232 = 8'he8 == io_addr[9:2] ? 32'h0 : _GEN_231; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_233 = 8'he9 == io_addr[9:2] ? 32'h0 : _GEN_232; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_234 = 8'hea == io_addr[9:2] ? 32'h0 : _GEN_233; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_235 = 8'heb == io_addr[9:2] ? 32'h0 : _GEN_234; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_236 = 8'hec == io_addr[9:2] ? 32'h0 : _GEN_235; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_237 = 8'hed == io_addr[9:2] ? 32'h0 : _GEN_236; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_238 = 8'hee == io_addr[9:2] ? 32'h0 : _GEN_237; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_239 = 8'hef == io_addr[9:2] ? 32'h0 : _GEN_238; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_240 = 8'hf0 == io_addr[9:2] ? 32'h0 : _GEN_239; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_241 = 8'hf1 == io_addr[9:2] ? 32'h0 : _GEN_240; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_242 = 8'hf2 == io_addr[9:2] ? 32'h0 : _GEN_241; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_243 = 8'hf3 == io_addr[9:2] ? 32'h0 : _GEN_242; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_244 = 8'hf4 == io_addr[9:2] ? 32'h0 : _GEN_243; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_245 = 8'hf5 == io_addr[9:2] ? 32'h0 : _GEN_244; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_246 = 8'hf6 == io_addr[9:2] ? 32'h0 : _GEN_245; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_247 = 8'hf7 == io_addr[9:2] ? 32'h0 : _GEN_246; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_248 = 8'hf8 == io_addr[9:2] ? 32'h0 : _GEN_247; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_249 = 8'hf9 == io_addr[9:2] ? 32'h0 : _GEN_248; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_250 = 8'hfa == io_addr[9:2] ? 32'h0 : _GEN_249; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_251 = 8'hfb == io_addr[9:2] ? 32'h0 : _GEN_250; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_252 = 8'hfc == io_addr[9:2] ? 32'h0 : _GEN_251; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_253 = 8'hfd == io_addr[9:2] ? 32'h0 : _GEN_252; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_254 = 8'hfe == io_addr[9:2] ? 32'h0 : _GEN_253; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_255 = 8'hff == io_addr[9:2] ? 32'h0 : _GEN_254; // @[InstMemory.scala 20:{11,11}]
  wire [8:0] _GEN_1024 = {{1'd0}, io_addr[9:2]}; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_256 = 9'h100 == _GEN_1024 ? 32'h0 : _GEN_255; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_257 = 9'h101 == _GEN_1024 ? 32'h0 : _GEN_256; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_258 = 9'h102 == _GEN_1024 ? 32'h0 : _GEN_257; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_259 = 9'h103 == _GEN_1024 ? 32'h0 : _GEN_258; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_260 = 9'h104 == _GEN_1024 ? 32'h0 : _GEN_259; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_261 = 9'h105 == _GEN_1024 ? 32'h0 : _GEN_260; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_262 = 9'h106 == _GEN_1024 ? 32'h0 : _GEN_261; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_263 = 9'h107 == _GEN_1024 ? 32'h0 : _GEN_262; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_264 = 9'h108 == _GEN_1024 ? 32'h0 : _GEN_263; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_265 = 9'h109 == _GEN_1024 ? 32'h0 : _GEN_264; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_266 = 9'h10a == _GEN_1024 ? 32'h0 : _GEN_265; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_267 = 9'h10b == _GEN_1024 ? 32'h0 : _GEN_266; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_268 = 9'h10c == _GEN_1024 ? 32'h0 : _GEN_267; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_269 = 9'h10d == _GEN_1024 ? 32'h0 : _GEN_268; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_270 = 9'h10e == _GEN_1024 ? 32'h0 : _GEN_269; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_271 = 9'h10f == _GEN_1024 ? 32'h0 : _GEN_270; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_272 = 9'h110 == _GEN_1024 ? 32'h0 : _GEN_271; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_273 = 9'h111 == _GEN_1024 ? 32'h0 : _GEN_272; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_274 = 9'h112 == _GEN_1024 ? 32'h0 : _GEN_273; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_275 = 9'h113 == _GEN_1024 ? 32'h0 : _GEN_274; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_276 = 9'h114 == _GEN_1024 ? 32'h0 : _GEN_275; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_277 = 9'h115 == _GEN_1024 ? 32'h0 : _GEN_276; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_278 = 9'h116 == _GEN_1024 ? 32'h0 : _GEN_277; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_279 = 9'h117 == _GEN_1024 ? 32'h0 : _GEN_278; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_280 = 9'h118 == _GEN_1024 ? 32'h0 : _GEN_279; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_281 = 9'h119 == _GEN_1024 ? 32'h0 : _GEN_280; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_282 = 9'h11a == _GEN_1024 ? 32'h0 : _GEN_281; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_283 = 9'h11b == _GEN_1024 ? 32'h0 : _GEN_282; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_284 = 9'h11c == _GEN_1024 ? 32'h0 : _GEN_283; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_285 = 9'h11d == _GEN_1024 ? 32'h0 : _GEN_284; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_286 = 9'h11e == _GEN_1024 ? 32'h0 : _GEN_285; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_287 = 9'h11f == _GEN_1024 ? 32'h0 : _GEN_286; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_288 = 9'h120 == _GEN_1024 ? 32'h0 : _GEN_287; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_289 = 9'h121 == _GEN_1024 ? 32'h0 : _GEN_288; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_290 = 9'h122 == _GEN_1024 ? 32'h0 : _GEN_289; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_291 = 9'h123 == _GEN_1024 ? 32'h0 : _GEN_290; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_292 = 9'h124 == _GEN_1024 ? 32'h0 : _GEN_291; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_293 = 9'h125 == _GEN_1024 ? 32'h0 : _GEN_292; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_294 = 9'h126 == _GEN_1024 ? 32'h0 : _GEN_293; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_295 = 9'h127 == _GEN_1024 ? 32'h0 : _GEN_294; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_296 = 9'h128 == _GEN_1024 ? 32'h0 : _GEN_295; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_297 = 9'h129 == _GEN_1024 ? 32'h0 : _GEN_296; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_298 = 9'h12a == _GEN_1024 ? 32'h0 : _GEN_297; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_299 = 9'h12b == _GEN_1024 ? 32'h0 : _GEN_298; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_300 = 9'h12c == _GEN_1024 ? 32'h0 : _GEN_299; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_301 = 9'h12d == _GEN_1024 ? 32'h0 : _GEN_300; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_302 = 9'h12e == _GEN_1024 ? 32'h0 : _GEN_301; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_303 = 9'h12f == _GEN_1024 ? 32'h0 : _GEN_302; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_304 = 9'h130 == _GEN_1024 ? 32'h0 : _GEN_303; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_305 = 9'h131 == _GEN_1024 ? 32'h0 : _GEN_304; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_306 = 9'h132 == _GEN_1024 ? 32'h0 : _GEN_305; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_307 = 9'h133 == _GEN_1024 ? 32'h0 : _GEN_306; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_308 = 9'h134 == _GEN_1024 ? 32'h0 : _GEN_307; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_309 = 9'h135 == _GEN_1024 ? 32'h0 : _GEN_308; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_310 = 9'h136 == _GEN_1024 ? 32'h0 : _GEN_309; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_311 = 9'h137 == _GEN_1024 ? 32'h0 : _GEN_310; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_312 = 9'h138 == _GEN_1024 ? 32'h0 : _GEN_311; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_313 = 9'h139 == _GEN_1024 ? 32'h0 : _GEN_312; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_314 = 9'h13a == _GEN_1024 ? 32'h0 : _GEN_313; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_315 = 9'h13b == _GEN_1024 ? 32'h0 : _GEN_314; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_316 = 9'h13c == _GEN_1024 ? 32'h0 : _GEN_315; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_317 = 9'h13d == _GEN_1024 ? 32'h0 : _GEN_316; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_318 = 9'h13e == _GEN_1024 ? 32'h0 : _GEN_317; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_319 = 9'h13f == _GEN_1024 ? 32'h0 : _GEN_318; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_320 = 9'h140 == _GEN_1024 ? 32'h0 : _GEN_319; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_321 = 9'h141 == _GEN_1024 ? 32'h0 : _GEN_320; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_322 = 9'h142 == _GEN_1024 ? 32'h0 : _GEN_321; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_323 = 9'h143 == _GEN_1024 ? 32'h0 : _GEN_322; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_324 = 9'h144 == _GEN_1024 ? 32'h0 : _GEN_323; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_325 = 9'h145 == _GEN_1024 ? 32'h0 : _GEN_324; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_326 = 9'h146 == _GEN_1024 ? 32'h0 : _GEN_325; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_327 = 9'h147 == _GEN_1024 ? 32'h0 : _GEN_326; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_328 = 9'h148 == _GEN_1024 ? 32'h0 : _GEN_327; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_329 = 9'h149 == _GEN_1024 ? 32'h0 : _GEN_328; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_330 = 9'h14a == _GEN_1024 ? 32'h0 : _GEN_329; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_331 = 9'h14b == _GEN_1024 ? 32'h0 : _GEN_330; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_332 = 9'h14c == _GEN_1024 ? 32'h0 : _GEN_331; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_333 = 9'h14d == _GEN_1024 ? 32'h0 : _GEN_332; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_334 = 9'h14e == _GEN_1024 ? 32'h0 : _GEN_333; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_335 = 9'h14f == _GEN_1024 ? 32'h0 : _GEN_334; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_336 = 9'h150 == _GEN_1024 ? 32'h0 : _GEN_335; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_337 = 9'h151 == _GEN_1024 ? 32'h0 : _GEN_336; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_338 = 9'h152 == _GEN_1024 ? 32'h0 : _GEN_337; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_339 = 9'h153 == _GEN_1024 ? 32'h0 : _GEN_338; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_340 = 9'h154 == _GEN_1024 ? 32'h0 : _GEN_339; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_341 = 9'h155 == _GEN_1024 ? 32'h0 : _GEN_340; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_342 = 9'h156 == _GEN_1024 ? 32'h0 : _GEN_341; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_343 = 9'h157 == _GEN_1024 ? 32'h0 : _GEN_342; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_344 = 9'h158 == _GEN_1024 ? 32'h0 : _GEN_343; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_345 = 9'h159 == _GEN_1024 ? 32'h0 : _GEN_344; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_346 = 9'h15a == _GEN_1024 ? 32'h0 : _GEN_345; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_347 = 9'h15b == _GEN_1024 ? 32'h0 : _GEN_346; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_348 = 9'h15c == _GEN_1024 ? 32'h0 : _GEN_347; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_349 = 9'h15d == _GEN_1024 ? 32'h0 : _GEN_348; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_350 = 9'h15e == _GEN_1024 ? 32'h0 : _GEN_349; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_351 = 9'h15f == _GEN_1024 ? 32'h0 : _GEN_350; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_352 = 9'h160 == _GEN_1024 ? 32'h0 : _GEN_351; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_353 = 9'h161 == _GEN_1024 ? 32'h0 : _GEN_352; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_354 = 9'h162 == _GEN_1024 ? 32'h0 : _GEN_353; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_355 = 9'h163 == _GEN_1024 ? 32'h0 : _GEN_354; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_356 = 9'h164 == _GEN_1024 ? 32'h0 : _GEN_355; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_357 = 9'h165 == _GEN_1024 ? 32'h0 : _GEN_356; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_358 = 9'h166 == _GEN_1024 ? 32'h0 : _GEN_357; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_359 = 9'h167 == _GEN_1024 ? 32'h0 : _GEN_358; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_360 = 9'h168 == _GEN_1024 ? 32'h0 : _GEN_359; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_361 = 9'h169 == _GEN_1024 ? 32'h0 : _GEN_360; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_362 = 9'h16a == _GEN_1024 ? 32'h0 : _GEN_361; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_363 = 9'h16b == _GEN_1024 ? 32'h0 : _GEN_362; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_364 = 9'h16c == _GEN_1024 ? 32'h0 : _GEN_363; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_365 = 9'h16d == _GEN_1024 ? 32'h0 : _GEN_364; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_366 = 9'h16e == _GEN_1024 ? 32'h0 : _GEN_365; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_367 = 9'h16f == _GEN_1024 ? 32'h0 : _GEN_366; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_368 = 9'h170 == _GEN_1024 ? 32'h0 : _GEN_367; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_369 = 9'h171 == _GEN_1024 ? 32'h0 : _GEN_368; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_370 = 9'h172 == _GEN_1024 ? 32'h0 : _GEN_369; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_371 = 9'h173 == _GEN_1024 ? 32'h0 : _GEN_370; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_372 = 9'h174 == _GEN_1024 ? 32'h0 : _GEN_371; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_373 = 9'h175 == _GEN_1024 ? 32'h0 : _GEN_372; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_374 = 9'h176 == _GEN_1024 ? 32'h0 : _GEN_373; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_375 = 9'h177 == _GEN_1024 ? 32'h0 : _GEN_374; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_376 = 9'h178 == _GEN_1024 ? 32'h0 : _GEN_375; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_377 = 9'h179 == _GEN_1024 ? 32'h0 : _GEN_376; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_378 = 9'h17a == _GEN_1024 ? 32'h0 : _GEN_377; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_379 = 9'h17b == _GEN_1024 ? 32'h0 : _GEN_378; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_380 = 9'h17c == _GEN_1024 ? 32'h0 : _GEN_379; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_381 = 9'h17d == _GEN_1024 ? 32'h0 : _GEN_380; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_382 = 9'h17e == _GEN_1024 ? 32'h0 : _GEN_381; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_383 = 9'h17f == _GEN_1024 ? 32'h0 : _GEN_382; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_384 = 9'h180 == _GEN_1024 ? 32'h0 : _GEN_383; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_385 = 9'h181 == _GEN_1024 ? 32'h0 : _GEN_384; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_386 = 9'h182 == _GEN_1024 ? 32'h0 : _GEN_385; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_387 = 9'h183 == _GEN_1024 ? 32'h0 : _GEN_386; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_388 = 9'h184 == _GEN_1024 ? 32'h0 : _GEN_387; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_389 = 9'h185 == _GEN_1024 ? 32'h0 : _GEN_388; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_390 = 9'h186 == _GEN_1024 ? 32'h0 : _GEN_389; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_391 = 9'h187 == _GEN_1024 ? 32'h0 : _GEN_390; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_392 = 9'h188 == _GEN_1024 ? 32'h0 : _GEN_391; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_393 = 9'h189 == _GEN_1024 ? 32'h0 : _GEN_392; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_394 = 9'h18a == _GEN_1024 ? 32'h0 : _GEN_393; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_395 = 9'h18b == _GEN_1024 ? 32'h0 : _GEN_394; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_396 = 9'h18c == _GEN_1024 ? 32'h0 : _GEN_395; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_397 = 9'h18d == _GEN_1024 ? 32'h0 : _GEN_396; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_398 = 9'h18e == _GEN_1024 ? 32'h0 : _GEN_397; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_399 = 9'h18f == _GEN_1024 ? 32'h0 : _GEN_398; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_400 = 9'h190 == _GEN_1024 ? 32'h0 : _GEN_399; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_401 = 9'h191 == _GEN_1024 ? 32'h0 : _GEN_400; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_402 = 9'h192 == _GEN_1024 ? 32'h0 : _GEN_401; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_403 = 9'h193 == _GEN_1024 ? 32'h0 : _GEN_402; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_404 = 9'h194 == _GEN_1024 ? 32'h0 : _GEN_403; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_405 = 9'h195 == _GEN_1024 ? 32'h0 : _GEN_404; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_406 = 9'h196 == _GEN_1024 ? 32'h0 : _GEN_405; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_407 = 9'h197 == _GEN_1024 ? 32'h0 : _GEN_406; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_408 = 9'h198 == _GEN_1024 ? 32'h0 : _GEN_407; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_409 = 9'h199 == _GEN_1024 ? 32'h0 : _GEN_408; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_410 = 9'h19a == _GEN_1024 ? 32'h0 : _GEN_409; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_411 = 9'h19b == _GEN_1024 ? 32'h0 : _GEN_410; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_412 = 9'h19c == _GEN_1024 ? 32'h0 : _GEN_411; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_413 = 9'h19d == _GEN_1024 ? 32'h0 : _GEN_412; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_414 = 9'h19e == _GEN_1024 ? 32'h0 : _GEN_413; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_415 = 9'h19f == _GEN_1024 ? 32'h0 : _GEN_414; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_416 = 9'h1a0 == _GEN_1024 ? 32'h0 : _GEN_415; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_417 = 9'h1a1 == _GEN_1024 ? 32'h0 : _GEN_416; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_418 = 9'h1a2 == _GEN_1024 ? 32'h0 : _GEN_417; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_419 = 9'h1a3 == _GEN_1024 ? 32'h0 : _GEN_418; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_420 = 9'h1a4 == _GEN_1024 ? 32'h0 : _GEN_419; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_421 = 9'h1a5 == _GEN_1024 ? 32'h0 : _GEN_420; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_422 = 9'h1a6 == _GEN_1024 ? 32'h0 : _GEN_421; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_423 = 9'h1a7 == _GEN_1024 ? 32'h0 : _GEN_422; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_424 = 9'h1a8 == _GEN_1024 ? 32'h0 : _GEN_423; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_425 = 9'h1a9 == _GEN_1024 ? 32'h0 : _GEN_424; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_426 = 9'h1aa == _GEN_1024 ? 32'h0 : _GEN_425; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_427 = 9'h1ab == _GEN_1024 ? 32'h0 : _GEN_426; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_428 = 9'h1ac == _GEN_1024 ? 32'h0 : _GEN_427; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_429 = 9'h1ad == _GEN_1024 ? 32'h0 : _GEN_428; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_430 = 9'h1ae == _GEN_1024 ? 32'h0 : _GEN_429; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_431 = 9'h1af == _GEN_1024 ? 32'h0 : _GEN_430; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_432 = 9'h1b0 == _GEN_1024 ? 32'h0 : _GEN_431; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_433 = 9'h1b1 == _GEN_1024 ? 32'h0 : _GEN_432; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_434 = 9'h1b2 == _GEN_1024 ? 32'h0 : _GEN_433; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_435 = 9'h1b3 == _GEN_1024 ? 32'h0 : _GEN_434; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_436 = 9'h1b4 == _GEN_1024 ? 32'h0 : _GEN_435; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_437 = 9'h1b5 == _GEN_1024 ? 32'h0 : _GEN_436; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_438 = 9'h1b6 == _GEN_1024 ? 32'h0 : _GEN_437; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_439 = 9'h1b7 == _GEN_1024 ? 32'h0 : _GEN_438; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_440 = 9'h1b8 == _GEN_1024 ? 32'h0 : _GEN_439; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_441 = 9'h1b9 == _GEN_1024 ? 32'h0 : _GEN_440; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_442 = 9'h1ba == _GEN_1024 ? 32'h0 : _GEN_441; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_443 = 9'h1bb == _GEN_1024 ? 32'h0 : _GEN_442; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_444 = 9'h1bc == _GEN_1024 ? 32'h0 : _GEN_443; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_445 = 9'h1bd == _GEN_1024 ? 32'h0 : _GEN_444; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_446 = 9'h1be == _GEN_1024 ? 32'h0 : _GEN_445; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_447 = 9'h1bf == _GEN_1024 ? 32'h0 : _GEN_446; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_448 = 9'h1c0 == _GEN_1024 ? 32'h0 : _GEN_447; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_449 = 9'h1c1 == _GEN_1024 ? 32'h0 : _GEN_448; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_450 = 9'h1c2 == _GEN_1024 ? 32'h0 : _GEN_449; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_451 = 9'h1c3 == _GEN_1024 ? 32'h0 : _GEN_450; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_452 = 9'h1c4 == _GEN_1024 ? 32'h0 : _GEN_451; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_453 = 9'h1c5 == _GEN_1024 ? 32'h0 : _GEN_452; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_454 = 9'h1c6 == _GEN_1024 ? 32'h0 : _GEN_453; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_455 = 9'h1c7 == _GEN_1024 ? 32'h0 : _GEN_454; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_456 = 9'h1c8 == _GEN_1024 ? 32'h0 : _GEN_455; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_457 = 9'h1c9 == _GEN_1024 ? 32'h0 : _GEN_456; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_458 = 9'h1ca == _GEN_1024 ? 32'h0 : _GEN_457; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_459 = 9'h1cb == _GEN_1024 ? 32'h0 : _GEN_458; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_460 = 9'h1cc == _GEN_1024 ? 32'h0 : _GEN_459; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_461 = 9'h1cd == _GEN_1024 ? 32'h0 : _GEN_460; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_462 = 9'h1ce == _GEN_1024 ? 32'h0 : _GEN_461; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_463 = 9'h1cf == _GEN_1024 ? 32'h0 : _GEN_462; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_464 = 9'h1d0 == _GEN_1024 ? 32'h0 : _GEN_463; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_465 = 9'h1d1 == _GEN_1024 ? 32'h0 : _GEN_464; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_466 = 9'h1d2 == _GEN_1024 ? 32'h0 : _GEN_465; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_467 = 9'h1d3 == _GEN_1024 ? 32'h0 : _GEN_466; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_468 = 9'h1d4 == _GEN_1024 ? 32'h0 : _GEN_467; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_469 = 9'h1d5 == _GEN_1024 ? 32'h0 : _GEN_468; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_470 = 9'h1d6 == _GEN_1024 ? 32'h0 : _GEN_469; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_471 = 9'h1d7 == _GEN_1024 ? 32'h0 : _GEN_470; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_472 = 9'h1d8 == _GEN_1024 ? 32'h0 : _GEN_471; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_473 = 9'h1d9 == _GEN_1024 ? 32'h0 : _GEN_472; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_474 = 9'h1da == _GEN_1024 ? 32'h0 : _GEN_473; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_475 = 9'h1db == _GEN_1024 ? 32'h0 : _GEN_474; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_476 = 9'h1dc == _GEN_1024 ? 32'h0 : _GEN_475; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_477 = 9'h1dd == _GEN_1024 ? 32'h0 : _GEN_476; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_478 = 9'h1de == _GEN_1024 ? 32'h0 : _GEN_477; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_479 = 9'h1df == _GEN_1024 ? 32'h0 : _GEN_478; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_480 = 9'h1e0 == _GEN_1024 ? 32'h0 : _GEN_479; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_481 = 9'h1e1 == _GEN_1024 ? 32'h0 : _GEN_480; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_482 = 9'h1e2 == _GEN_1024 ? 32'h0 : _GEN_481; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_483 = 9'h1e3 == _GEN_1024 ? 32'h0 : _GEN_482; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_484 = 9'h1e4 == _GEN_1024 ? 32'h0 : _GEN_483; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_485 = 9'h1e5 == _GEN_1024 ? 32'h0 : _GEN_484; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_486 = 9'h1e6 == _GEN_1024 ? 32'h0 : _GEN_485; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_487 = 9'h1e7 == _GEN_1024 ? 32'h0 : _GEN_486; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_488 = 9'h1e8 == _GEN_1024 ? 32'h0 : _GEN_487; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_489 = 9'h1e9 == _GEN_1024 ? 32'h0 : _GEN_488; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_490 = 9'h1ea == _GEN_1024 ? 32'h0 : _GEN_489; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_491 = 9'h1eb == _GEN_1024 ? 32'h0 : _GEN_490; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_492 = 9'h1ec == _GEN_1024 ? 32'h0 : _GEN_491; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_493 = 9'h1ed == _GEN_1024 ? 32'h0 : _GEN_492; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_494 = 9'h1ee == _GEN_1024 ? 32'h0 : _GEN_493; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_495 = 9'h1ef == _GEN_1024 ? 32'h0 : _GEN_494; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_496 = 9'h1f0 == _GEN_1024 ? 32'h0 : _GEN_495; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_497 = 9'h1f1 == _GEN_1024 ? 32'h0 : _GEN_496; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_498 = 9'h1f2 == _GEN_1024 ? 32'h0 : _GEN_497; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_499 = 9'h1f3 == _GEN_1024 ? 32'h0 : _GEN_498; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_500 = 9'h1f4 == _GEN_1024 ? 32'h0 : _GEN_499; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_501 = 9'h1f5 == _GEN_1024 ? 32'h0 : _GEN_500; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_502 = 9'h1f6 == _GEN_1024 ? 32'h0 : _GEN_501; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_503 = 9'h1f7 == _GEN_1024 ? 32'h0 : _GEN_502; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_504 = 9'h1f8 == _GEN_1024 ? 32'h0 : _GEN_503; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_505 = 9'h1f9 == _GEN_1024 ? 32'h0 : _GEN_504; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_506 = 9'h1fa == _GEN_1024 ? 32'h0 : _GEN_505; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_507 = 9'h1fb == _GEN_1024 ? 32'h0 : _GEN_506; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_508 = 9'h1fc == _GEN_1024 ? 32'h0 : _GEN_507; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_509 = 9'h1fd == _GEN_1024 ? 32'h0 : _GEN_508; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_510 = 9'h1fe == _GEN_1024 ? 32'h0 : _GEN_509; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_511 = 9'h1ff == _GEN_1024 ? 32'h0 : _GEN_510; // @[InstMemory.scala 20:{11,11}]
  wire [9:0] _GEN_1280 = {{2'd0}, io_addr[9:2]}; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_512 = 10'h200 == _GEN_1280 ? 32'h0 : _GEN_511; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_513 = 10'h201 == _GEN_1280 ? 32'h0 : _GEN_512; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_514 = 10'h202 == _GEN_1280 ? 32'h0 : _GEN_513; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_515 = 10'h203 == _GEN_1280 ? 32'h0 : _GEN_514; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_516 = 10'h204 == _GEN_1280 ? 32'h0 : _GEN_515; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_517 = 10'h205 == _GEN_1280 ? 32'h0 : _GEN_516; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_518 = 10'h206 == _GEN_1280 ? 32'h0 : _GEN_517; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_519 = 10'h207 == _GEN_1280 ? 32'h0 : _GEN_518; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_520 = 10'h208 == _GEN_1280 ? 32'h0 : _GEN_519; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_521 = 10'h209 == _GEN_1280 ? 32'h0 : _GEN_520; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_522 = 10'h20a == _GEN_1280 ? 32'h0 : _GEN_521; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_523 = 10'h20b == _GEN_1280 ? 32'h0 : _GEN_522; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_524 = 10'h20c == _GEN_1280 ? 32'h0 : _GEN_523; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_525 = 10'h20d == _GEN_1280 ? 32'h0 : _GEN_524; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_526 = 10'h20e == _GEN_1280 ? 32'h0 : _GEN_525; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_527 = 10'h20f == _GEN_1280 ? 32'h0 : _GEN_526; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_528 = 10'h210 == _GEN_1280 ? 32'h0 : _GEN_527; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_529 = 10'h211 == _GEN_1280 ? 32'h0 : _GEN_528; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_530 = 10'h212 == _GEN_1280 ? 32'h0 : _GEN_529; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_531 = 10'h213 == _GEN_1280 ? 32'h0 : _GEN_530; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_532 = 10'h214 == _GEN_1280 ? 32'h0 : _GEN_531; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_533 = 10'h215 == _GEN_1280 ? 32'h0 : _GEN_532; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_534 = 10'h216 == _GEN_1280 ? 32'h0 : _GEN_533; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_535 = 10'h217 == _GEN_1280 ? 32'h0 : _GEN_534; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_536 = 10'h218 == _GEN_1280 ? 32'h0 : _GEN_535; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_537 = 10'h219 == _GEN_1280 ? 32'h0 : _GEN_536; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_538 = 10'h21a == _GEN_1280 ? 32'h0 : _GEN_537; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_539 = 10'h21b == _GEN_1280 ? 32'h0 : _GEN_538; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_540 = 10'h21c == _GEN_1280 ? 32'h0 : _GEN_539; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_541 = 10'h21d == _GEN_1280 ? 32'h0 : _GEN_540; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_542 = 10'h21e == _GEN_1280 ? 32'h0 : _GEN_541; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_543 = 10'h21f == _GEN_1280 ? 32'h0 : _GEN_542; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_544 = 10'h220 == _GEN_1280 ? 32'h0 : _GEN_543; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_545 = 10'h221 == _GEN_1280 ? 32'h0 : _GEN_544; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_546 = 10'h222 == _GEN_1280 ? 32'h0 : _GEN_545; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_547 = 10'h223 == _GEN_1280 ? 32'h0 : _GEN_546; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_548 = 10'h224 == _GEN_1280 ? 32'h0 : _GEN_547; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_549 = 10'h225 == _GEN_1280 ? 32'h0 : _GEN_548; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_550 = 10'h226 == _GEN_1280 ? 32'h0 : _GEN_549; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_551 = 10'h227 == _GEN_1280 ? 32'h0 : _GEN_550; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_552 = 10'h228 == _GEN_1280 ? 32'h0 : _GEN_551; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_553 = 10'h229 == _GEN_1280 ? 32'h0 : _GEN_552; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_554 = 10'h22a == _GEN_1280 ? 32'h0 : _GEN_553; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_555 = 10'h22b == _GEN_1280 ? 32'h0 : _GEN_554; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_556 = 10'h22c == _GEN_1280 ? 32'h0 : _GEN_555; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_557 = 10'h22d == _GEN_1280 ? 32'h0 : _GEN_556; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_558 = 10'h22e == _GEN_1280 ? 32'h0 : _GEN_557; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_559 = 10'h22f == _GEN_1280 ? 32'h0 : _GEN_558; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_560 = 10'h230 == _GEN_1280 ? 32'h0 : _GEN_559; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_561 = 10'h231 == _GEN_1280 ? 32'h0 : _GEN_560; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_562 = 10'h232 == _GEN_1280 ? 32'h0 : _GEN_561; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_563 = 10'h233 == _GEN_1280 ? 32'h0 : _GEN_562; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_564 = 10'h234 == _GEN_1280 ? 32'h0 : _GEN_563; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_565 = 10'h235 == _GEN_1280 ? 32'h0 : _GEN_564; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_566 = 10'h236 == _GEN_1280 ? 32'h0 : _GEN_565; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_567 = 10'h237 == _GEN_1280 ? 32'h0 : _GEN_566; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_568 = 10'h238 == _GEN_1280 ? 32'h0 : _GEN_567; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_569 = 10'h239 == _GEN_1280 ? 32'h0 : _GEN_568; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_570 = 10'h23a == _GEN_1280 ? 32'h0 : _GEN_569; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_571 = 10'h23b == _GEN_1280 ? 32'h0 : _GEN_570; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_572 = 10'h23c == _GEN_1280 ? 32'h0 : _GEN_571; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_573 = 10'h23d == _GEN_1280 ? 32'h0 : _GEN_572; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_574 = 10'h23e == _GEN_1280 ? 32'h0 : _GEN_573; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_575 = 10'h23f == _GEN_1280 ? 32'h0 : _GEN_574; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_576 = 10'h240 == _GEN_1280 ? 32'h0 : _GEN_575; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_577 = 10'h241 == _GEN_1280 ? 32'h0 : _GEN_576; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_578 = 10'h242 == _GEN_1280 ? 32'h0 : _GEN_577; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_579 = 10'h243 == _GEN_1280 ? 32'h0 : _GEN_578; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_580 = 10'h244 == _GEN_1280 ? 32'h0 : _GEN_579; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_581 = 10'h245 == _GEN_1280 ? 32'h0 : _GEN_580; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_582 = 10'h246 == _GEN_1280 ? 32'h0 : _GEN_581; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_583 = 10'h247 == _GEN_1280 ? 32'h0 : _GEN_582; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_584 = 10'h248 == _GEN_1280 ? 32'h0 : _GEN_583; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_585 = 10'h249 == _GEN_1280 ? 32'h0 : _GEN_584; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_586 = 10'h24a == _GEN_1280 ? 32'h0 : _GEN_585; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_587 = 10'h24b == _GEN_1280 ? 32'h0 : _GEN_586; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_588 = 10'h24c == _GEN_1280 ? 32'h0 : _GEN_587; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_589 = 10'h24d == _GEN_1280 ? 32'h0 : _GEN_588; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_590 = 10'h24e == _GEN_1280 ? 32'h0 : _GEN_589; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_591 = 10'h24f == _GEN_1280 ? 32'h0 : _GEN_590; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_592 = 10'h250 == _GEN_1280 ? 32'h0 : _GEN_591; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_593 = 10'h251 == _GEN_1280 ? 32'h0 : _GEN_592; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_594 = 10'h252 == _GEN_1280 ? 32'h0 : _GEN_593; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_595 = 10'h253 == _GEN_1280 ? 32'h0 : _GEN_594; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_596 = 10'h254 == _GEN_1280 ? 32'h0 : _GEN_595; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_597 = 10'h255 == _GEN_1280 ? 32'h0 : _GEN_596; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_598 = 10'h256 == _GEN_1280 ? 32'h0 : _GEN_597; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_599 = 10'h257 == _GEN_1280 ? 32'h0 : _GEN_598; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_600 = 10'h258 == _GEN_1280 ? 32'h0 : _GEN_599; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_601 = 10'h259 == _GEN_1280 ? 32'h0 : _GEN_600; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_602 = 10'h25a == _GEN_1280 ? 32'h0 : _GEN_601; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_603 = 10'h25b == _GEN_1280 ? 32'h0 : _GEN_602; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_604 = 10'h25c == _GEN_1280 ? 32'h0 : _GEN_603; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_605 = 10'h25d == _GEN_1280 ? 32'h0 : _GEN_604; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_606 = 10'h25e == _GEN_1280 ? 32'h0 : _GEN_605; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_607 = 10'h25f == _GEN_1280 ? 32'h0 : _GEN_606; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_608 = 10'h260 == _GEN_1280 ? 32'h0 : _GEN_607; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_609 = 10'h261 == _GEN_1280 ? 32'h0 : _GEN_608; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_610 = 10'h262 == _GEN_1280 ? 32'h0 : _GEN_609; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_611 = 10'h263 == _GEN_1280 ? 32'h0 : _GEN_610; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_612 = 10'h264 == _GEN_1280 ? 32'h0 : _GEN_611; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_613 = 10'h265 == _GEN_1280 ? 32'h0 : _GEN_612; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_614 = 10'h266 == _GEN_1280 ? 32'h0 : _GEN_613; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_615 = 10'h267 == _GEN_1280 ? 32'h0 : _GEN_614; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_616 = 10'h268 == _GEN_1280 ? 32'h0 : _GEN_615; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_617 = 10'h269 == _GEN_1280 ? 32'h0 : _GEN_616; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_618 = 10'h26a == _GEN_1280 ? 32'h0 : _GEN_617; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_619 = 10'h26b == _GEN_1280 ? 32'h0 : _GEN_618; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_620 = 10'h26c == _GEN_1280 ? 32'h0 : _GEN_619; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_621 = 10'h26d == _GEN_1280 ? 32'h0 : _GEN_620; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_622 = 10'h26e == _GEN_1280 ? 32'h0 : _GEN_621; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_623 = 10'h26f == _GEN_1280 ? 32'h0 : _GEN_622; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_624 = 10'h270 == _GEN_1280 ? 32'h0 : _GEN_623; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_625 = 10'h271 == _GEN_1280 ? 32'h0 : _GEN_624; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_626 = 10'h272 == _GEN_1280 ? 32'h0 : _GEN_625; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_627 = 10'h273 == _GEN_1280 ? 32'h0 : _GEN_626; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_628 = 10'h274 == _GEN_1280 ? 32'h0 : _GEN_627; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_629 = 10'h275 == _GEN_1280 ? 32'h0 : _GEN_628; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_630 = 10'h276 == _GEN_1280 ? 32'h0 : _GEN_629; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_631 = 10'h277 == _GEN_1280 ? 32'h0 : _GEN_630; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_632 = 10'h278 == _GEN_1280 ? 32'h0 : _GEN_631; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_633 = 10'h279 == _GEN_1280 ? 32'h0 : _GEN_632; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_634 = 10'h27a == _GEN_1280 ? 32'h0 : _GEN_633; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_635 = 10'h27b == _GEN_1280 ? 32'h0 : _GEN_634; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_636 = 10'h27c == _GEN_1280 ? 32'h0 : _GEN_635; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_637 = 10'h27d == _GEN_1280 ? 32'h0 : _GEN_636; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_638 = 10'h27e == _GEN_1280 ? 32'h0 : _GEN_637; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_639 = 10'h27f == _GEN_1280 ? 32'h0 : _GEN_638; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_640 = 10'h280 == _GEN_1280 ? 32'h0 : _GEN_639; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_641 = 10'h281 == _GEN_1280 ? 32'h0 : _GEN_640; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_642 = 10'h282 == _GEN_1280 ? 32'h0 : _GEN_641; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_643 = 10'h283 == _GEN_1280 ? 32'h0 : _GEN_642; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_644 = 10'h284 == _GEN_1280 ? 32'h0 : _GEN_643; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_645 = 10'h285 == _GEN_1280 ? 32'h0 : _GEN_644; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_646 = 10'h286 == _GEN_1280 ? 32'h0 : _GEN_645; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_647 = 10'h287 == _GEN_1280 ? 32'h0 : _GEN_646; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_648 = 10'h288 == _GEN_1280 ? 32'h0 : _GEN_647; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_649 = 10'h289 == _GEN_1280 ? 32'h0 : _GEN_648; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_650 = 10'h28a == _GEN_1280 ? 32'h0 : _GEN_649; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_651 = 10'h28b == _GEN_1280 ? 32'h0 : _GEN_650; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_652 = 10'h28c == _GEN_1280 ? 32'h0 : _GEN_651; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_653 = 10'h28d == _GEN_1280 ? 32'h0 : _GEN_652; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_654 = 10'h28e == _GEN_1280 ? 32'h0 : _GEN_653; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_655 = 10'h28f == _GEN_1280 ? 32'h0 : _GEN_654; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_656 = 10'h290 == _GEN_1280 ? 32'h0 : _GEN_655; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_657 = 10'h291 == _GEN_1280 ? 32'h0 : _GEN_656; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_658 = 10'h292 == _GEN_1280 ? 32'h0 : _GEN_657; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_659 = 10'h293 == _GEN_1280 ? 32'h0 : _GEN_658; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_660 = 10'h294 == _GEN_1280 ? 32'h0 : _GEN_659; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_661 = 10'h295 == _GEN_1280 ? 32'h0 : _GEN_660; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_662 = 10'h296 == _GEN_1280 ? 32'h0 : _GEN_661; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_663 = 10'h297 == _GEN_1280 ? 32'h0 : _GEN_662; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_664 = 10'h298 == _GEN_1280 ? 32'h0 : _GEN_663; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_665 = 10'h299 == _GEN_1280 ? 32'h0 : _GEN_664; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_666 = 10'h29a == _GEN_1280 ? 32'h0 : _GEN_665; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_667 = 10'h29b == _GEN_1280 ? 32'h0 : _GEN_666; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_668 = 10'h29c == _GEN_1280 ? 32'h0 : _GEN_667; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_669 = 10'h29d == _GEN_1280 ? 32'h0 : _GEN_668; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_670 = 10'h29e == _GEN_1280 ? 32'h0 : _GEN_669; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_671 = 10'h29f == _GEN_1280 ? 32'h0 : _GEN_670; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_672 = 10'h2a0 == _GEN_1280 ? 32'h0 : _GEN_671; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_673 = 10'h2a1 == _GEN_1280 ? 32'h0 : _GEN_672; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_674 = 10'h2a2 == _GEN_1280 ? 32'h0 : _GEN_673; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_675 = 10'h2a3 == _GEN_1280 ? 32'h0 : _GEN_674; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_676 = 10'h2a4 == _GEN_1280 ? 32'h0 : _GEN_675; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_677 = 10'h2a5 == _GEN_1280 ? 32'h0 : _GEN_676; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_678 = 10'h2a6 == _GEN_1280 ? 32'h0 : _GEN_677; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_679 = 10'h2a7 == _GEN_1280 ? 32'h0 : _GEN_678; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_680 = 10'h2a8 == _GEN_1280 ? 32'h0 : _GEN_679; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_681 = 10'h2a9 == _GEN_1280 ? 32'h0 : _GEN_680; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_682 = 10'h2aa == _GEN_1280 ? 32'h0 : _GEN_681; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_683 = 10'h2ab == _GEN_1280 ? 32'h0 : _GEN_682; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_684 = 10'h2ac == _GEN_1280 ? 32'h0 : _GEN_683; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_685 = 10'h2ad == _GEN_1280 ? 32'h0 : _GEN_684; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_686 = 10'h2ae == _GEN_1280 ? 32'h0 : _GEN_685; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_687 = 10'h2af == _GEN_1280 ? 32'h0 : _GEN_686; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_688 = 10'h2b0 == _GEN_1280 ? 32'h0 : _GEN_687; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_689 = 10'h2b1 == _GEN_1280 ? 32'h0 : _GEN_688; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_690 = 10'h2b2 == _GEN_1280 ? 32'h0 : _GEN_689; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_691 = 10'h2b3 == _GEN_1280 ? 32'h0 : _GEN_690; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_692 = 10'h2b4 == _GEN_1280 ? 32'h0 : _GEN_691; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_693 = 10'h2b5 == _GEN_1280 ? 32'h0 : _GEN_692; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_694 = 10'h2b6 == _GEN_1280 ? 32'h0 : _GEN_693; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_695 = 10'h2b7 == _GEN_1280 ? 32'h0 : _GEN_694; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_696 = 10'h2b8 == _GEN_1280 ? 32'h0 : _GEN_695; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_697 = 10'h2b9 == _GEN_1280 ? 32'h0 : _GEN_696; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_698 = 10'h2ba == _GEN_1280 ? 32'h0 : _GEN_697; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_699 = 10'h2bb == _GEN_1280 ? 32'h0 : _GEN_698; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_700 = 10'h2bc == _GEN_1280 ? 32'h0 : _GEN_699; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_701 = 10'h2bd == _GEN_1280 ? 32'h0 : _GEN_700; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_702 = 10'h2be == _GEN_1280 ? 32'h0 : _GEN_701; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_703 = 10'h2bf == _GEN_1280 ? 32'h0 : _GEN_702; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_704 = 10'h2c0 == _GEN_1280 ? 32'h0 : _GEN_703; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_705 = 10'h2c1 == _GEN_1280 ? 32'h0 : _GEN_704; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_706 = 10'h2c2 == _GEN_1280 ? 32'h0 : _GEN_705; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_707 = 10'h2c3 == _GEN_1280 ? 32'h0 : _GEN_706; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_708 = 10'h2c4 == _GEN_1280 ? 32'h0 : _GEN_707; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_709 = 10'h2c5 == _GEN_1280 ? 32'h0 : _GEN_708; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_710 = 10'h2c6 == _GEN_1280 ? 32'h0 : _GEN_709; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_711 = 10'h2c7 == _GEN_1280 ? 32'h0 : _GEN_710; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_712 = 10'h2c8 == _GEN_1280 ? 32'h0 : _GEN_711; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_713 = 10'h2c9 == _GEN_1280 ? 32'h0 : _GEN_712; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_714 = 10'h2ca == _GEN_1280 ? 32'h0 : _GEN_713; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_715 = 10'h2cb == _GEN_1280 ? 32'h0 : _GEN_714; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_716 = 10'h2cc == _GEN_1280 ? 32'h0 : _GEN_715; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_717 = 10'h2cd == _GEN_1280 ? 32'h0 : _GEN_716; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_718 = 10'h2ce == _GEN_1280 ? 32'h0 : _GEN_717; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_719 = 10'h2cf == _GEN_1280 ? 32'h0 : _GEN_718; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_720 = 10'h2d0 == _GEN_1280 ? 32'h0 : _GEN_719; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_721 = 10'h2d1 == _GEN_1280 ? 32'h0 : _GEN_720; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_722 = 10'h2d2 == _GEN_1280 ? 32'h0 : _GEN_721; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_723 = 10'h2d3 == _GEN_1280 ? 32'h0 : _GEN_722; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_724 = 10'h2d4 == _GEN_1280 ? 32'h0 : _GEN_723; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_725 = 10'h2d5 == _GEN_1280 ? 32'h0 : _GEN_724; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_726 = 10'h2d6 == _GEN_1280 ? 32'h0 : _GEN_725; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_727 = 10'h2d7 == _GEN_1280 ? 32'h0 : _GEN_726; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_728 = 10'h2d8 == _GEN_1280 ? 32'h0 : _GEN_727; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_729 = 10'h2d9 == _GEN_1280 ? 32'h0 : _GEN_728; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_730 = 10'h2da == _GEN_1280 ? 32'h0 : _GEN_729; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_731 = 10'h2db == _GEN_1280 ? 32'h0 : _GEN_730; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_732 = 10'h2dc == _GEN_1280 ? 32'h0 : _GEN_731; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_733 = 10'h2dd == _GEN_1280 ? 32'h0 : _GEN_732; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_734 = 10'h2de == _GEN_1280 ? 32'h0 : _GEN_733; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_735 = 10'h2df == _GEN_1280 ? 32'h0 : _GEN_734; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_736 = 10'h2e0 == _GEN_1280 ? 32'h0 : _GEN_735; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_737 = 10'h2e1 == _GEN_1280 ? 32'h0 : _GEN_736; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_738 = 10'h2e2 == _GEN_1280 ? 32'h0 : _GEN_737; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_739 = 10'h2e3 == _GEN_1280 ? 32'h0 : _GEN_738; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_740 = 10'h2e4 == _GEN_1280 ? 32'h0 : _GEN_739; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_741 = 10'h2e5 == _GEN_1280 ? 32'h0 : _GEN_740; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_742 = 10'h2e6 == _GEN_1280 ? 32'h0 : _GEN_741; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_743 = 10'h2e7 == _GEN_1280 ? 32'h0 : _GEN_742; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_744 = 10'h2e8 == _GEN_1280 ? 32'h0 : _GEN_743; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_745 = 10'h2e9 == _GEN_1280 ? 32'h0 : _GEN_744; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_746 = 10'h2ea == _GEN_1280 ? 32'h0 : _GEN_745; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_747 = 10'h2eb == _GEN_1280 ? 32'h0 : _GEN_746; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_748 = 10'h2ec == _GEN_1280 ? 32'h0 : _GEN_747; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_749 = 10'h2ed == _GEN_1280 ? 32'h0 : _GEN_748; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_750 = 10'h2ee == _GEN_1280 ? 32'h0 : _GEN_749; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_751 = 10'h2ef == _GEN_1280 ? 32'h0 : _GEN_750; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_752 = 10'h2f0 == _GEN_1280 ? 32'h0 : _GEN_751; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_753 = 10'h2f1 == _GEN_1280 ? 32'h0 : _GEN_752; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_754 = 10'h2f2 == _GEN_1280 ? 32'h0 : _GEN_753; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_755 = 10'h2f3 == _GEN_1280 ? 32'h0 : _GEN_754; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_756 = 10'h2f4 == _GEN_1280 ? 32'h0 : _GEN_755; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_757 = 10'h2f5 == _GEN_1280 ? 32'h0 : _GEN_756; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_758 = 10'h2f6 == _GEN_1280 ? 32'h0 : _GEN_757; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_759 = 10'h2f7 == _GEN_1280 ? 32'h0 : _GEN_758; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_760 = 10'h2f8 == _GEN_1280 ? 32'h0 : _GEN_759; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_761 = 10'h2f9 == _GEN_1280 ? 32'h0 : _GEN_760; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_762 = 10'h2fa == _GEN_1280 ? 32'h0 : _GEN_761; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_763 = 10'h2fb == _GEN_1280 ? 32'h0 : _GEN_762; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_764 = 10'h2fc == _GEN_1280 ? 32'h0 : _GEN_763; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_765 = 10'h2fd == _GEN_1280 ? 32'h0 : _GEN_764; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_766 = 10'h2fe == _GEN_1280 ? 32'h0 : _GEN_765; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_767 = 10'h2ff == _GEN_1280 ? 32'h0 : _GEN_766; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_768 = 10'h300 == _GEN_1280 ? 32'h0 : _GEN_767; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_769 = 10'h301 == _GEN_1280 ? 32'h0 : _GEN_768; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_770 = 10'h302 == _GEN_1280 ? 32'h0 : _GEN_769; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_771 = 10'h303 == _GEN_1280 ? 32'h0 : _GEN_770; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_772 = 10'h304 == _GEN_1280 ? 32'h0 : _GEN_771; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_773 = 10'h305 == _GEN_1280 ? 32'h0 : _GEN_772; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_774 = 10'h306 == _GEN_1280 ? 32'h0 : _GEN_773; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_775 = 10'h307 == _GEN_1280 ? 32'h0 : _GEN_774; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_776 = 10'h308 == _GEN_1280 ? 32'h0 : _GEN_775; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_777 = 10'h309 == _GEN_1280 ? 32'h0 : _GEN_776; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_778 = 10'h30a == _GEN_1280 ? 32'h0 : _GEN_777; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_779 = 10'h30b == _GEN_1280 ? 32'h0 : _GEN_778; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_780 = 10'h30c == _GEN_1280 ? 32'h0 : _GEN_779; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_781 = 10'h30d == _GEN_1280 ? 32'h0 : _GEN_780; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_782 = 10'h30e == _GEN_1280 ? 32'h0 : _GEN_781; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_783 = 10'h30f == _GEN_1280 ? 32'h0 : _GEN_782; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_784 = 10'h310 == _GEN_1280 ? 32'h0 : _GEN_783; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_785 = 10'h311 == _GEN_1280 ? 32'h0 : _GEN_784; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_786 = 10'h312 == _GEN_1280 ? 32'h0 : _GEN_785; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_787 = 10'h313 == _GEN_1280 ? 32'h0 : _GEN_786; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_788 = 10'h314 == _GEN_1280 ? 32'h0 : _GEN_787; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_789 = 10'h315 == _GEN_1280 ? 32'h0 : _GEN_788; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_790 = 10'h316 == _GEN_1280 ? 32'h0 : _GEN_789; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_791 = 10'h317 == _GEN_1280 ? 32'h0 : _GEN_790; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_792 = 10'h318 == _GEN_1280 ? 32'h0 : _GEN_791; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_793 = 10'h319 == _GEN_1280 ? 32'h0 : _GEN_792; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_794 = 10'h31a == _GEN_1280 ? 32'h0 : _GEN_793; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_795 = 10'h31b == _GEN_1280 ? 32'h0 : _GEN_794; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_796 = 10'h31c == _GEN_1280 ? 32'h0 : _GEN_795; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_797 = 10'h31d == _GEN_1280 ? 32'h0 : _GEN_796; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_798 = 10'h31e == _GEN_1280 ? 32'h0 : _GEN_797; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_799 = 10'h31f == _GEN_1280 ? 32'h0 : _GEN_798; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_800 = 10'h320 == _GEN_1280 ? 32'h0 : _GEN_799; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_801 = 10'h321 == _GEN_1280 ? 32'h0 : _GEN_800; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_802 = 10'h322 == _GEN_1280 ? 32'h0 : _GEN_801; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_803 = 10'h323 == _GEN_1280 ? 32'h0 : _GEN_802; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_804 = 10'h324 == _GEN_1280 ? 32'h0 : _GEN_803; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_805 = 10'h325 == _GEN_1280 ? 32'h0 : _GEN_804; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_806 = 10'h326 == _GEN_1280 ? 32'h0 : _GEN_805; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_807 = 10'h327 == _GEN_1280 ? 32'h0 : _GEN_806; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_808 = 10'h328 == _GEN_1280 ? 32'h0 : _GEN_807; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_809 = 10'h329 == _GEN_1280 ? 32'h0 : _GEN_808; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_810 = 10'h32a == _GEN_1280 ? 32'h0 : _GEN_809; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_811 = 10'h32b == _GEN_1280 ? 32'h0 : _GEN_810; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_812 = 10'h32c == _GEN_1280 ? 32'h0 : _GEN_811; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_813 = 10'h32d == _GEN_1280 ? 32'h0 : _GEN_812; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_814 = 10'h32e == _GEN_1280 ? 32'h0 : _GEN_813; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_815 = 10'h32f == _GEN_1280 ? 32'h0 : _GEN_814; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_816 = 10'h330 == _GEN_1280 ? 32'h0 : _GEN_815; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_817 = 10'h331 == _GEN_1280 ? 32'h0 : _GEN_816; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_818 = 10'h332 == _GEN_1280 ? 32'h0 : _GEN_817; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_819 = 10'h333 == _GEN_1280 ? 32'h0 : _GEN_818; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_820 = 10'h334 == _GEN_1280 ? 32'h0 : _GEN_819; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_821 = 10'h335 == _GEN_1280 ? 32'h0 : _GEN_820; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_822 = 10'h336 == _GEN_1280 ? 32'h0 : _GEN_821; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_823 = 10'h337 == _GEN_1280 ? 32'h0 : _GEN_822; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_824 = 10'h338 == _GEN_1280 ? 32'h0 : _GEN_823; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_825 = 10'h339 == _GEN_1280 ? 32'h0 : _GEN_824; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_826 = 10'h33a == _GEN_1280 ? 32'h0 : _GEN_825; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_827 = 10'h33b == _GEN_1280 ? 32'h0 : _GEN_826; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_828 = 10'h33c == _GEN_1280 ? 32'h0 : _GEN_827; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_829 = 10'h33d == _GEN_1280 ? 32'h0 : _GEN_828; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_830 = 10'h33e == _GEN_1280 ? 32'h0 : _GEN_829; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_831 = 10'h33f == _GEN_1280 ? 32'h0 : _GEN_830; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_832 = 10'h340 == _GEN_1280 ? 32'h0 : _GEN_831; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_833 = 10'h341 == _GEN_1280 ? 32'h0 : _GEN_832; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_834 = 10'h342 == _GEN_1280 ? 32'h0 : _GEN_833; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_835 = 10'h343 == _GEN_1280 ? 32'h0 : _GEN_834; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_836 = 10'h344 == _GEN_1280 ? 32'h0 : _GEN_835; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_837 = 10'h345 == _GEN_1280 ? 32'h0 : _GEN_836; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_838 = 10'h346 == _GEN_1280 ? 32'h0 : _GEN_837; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_839 = 10'h347 == _GEN_1280 ? 32'h0 : _GEN_838; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_840 = 10'h348 == _GEN_1280 ? 32'h0 : _GEN_839; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_841 = 10'h349 == _GEN_1280 ? 32'h0 : _GEN_840; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_842 = 10'h34a == _GEN_1280 ? 32'h0 : _GEN_841; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_843 = 10'h34b == _GEN_1280 ? 32'h0 : _GEN_842; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_844 = 10'h34c == _GEN_1280 ? 32'h0 : _GEN_843; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_845 = 10'h34d == _GEN_1280 ? 32'h0 : _GEN_844; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_846 = 10'h34e == _GEN_1280 ? 32'h0 : _GEN_845; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_847 = 10'h34f == _GEN_1280 ? 32'h0 : _GEN_846; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_848 = 10'h350 == _GEN_1280 ? 32'h0 : _GEN_847; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_849 = 10'h351 == _GEN_1280 ? 32'h0 : _GEN_848; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_850 = 10'h352 == _GEN_1280 ? 32'h0 : _GEN_849; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_851 = 10'h353 == _GEN_1280 ? 32'h0 : _GEN_850; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_852 = 10'h354 == _GEN_1280 ? 32'h0 : _GEN_851; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_853 = 10'h355 == _GEN_1280 ? 32'h0 : _GEN_852; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_854 = 10'h356 == _GEN_1280 ? 32'h0 : _GEN_853; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_855 = 10'h357 == _GEN_1280 ? 32'h0 : _GEN_854; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_856 = 10'h358 == _GEN_1280 ? 32'h0 : _GEN_855; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_857 = 10'h359 == _GEN_1280 ? 32'h0 : _GEN_856; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_858 = 10'h35a == _GEN_1280 ? 32'h0 : _GEN_857; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_859 = 10'h35b == _GEN_1280 ? 32'h0 : _GEN_858; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_860 = 10'h35c == _GEN_1280 ? 32'h0 : _GEN_859; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_861 = 10'h35d == _GEN_1280 ? 32'h0 : _GEN_860; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_862 = 10'h35e == _GEN_1280 ? 32'h0 : _GEN_861; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_863 = 10'h35f == _GEN_1280 ? 32'h0 : _GEN_862; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_864 = 10'h360 == _GEN_1280 ? 32'h0 : _GEN_863; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_865 = 10'h361 == _GEN_1280 ? 32'h0 : _GEN_864; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_866 = 10'h362 == _GEN_1280 ? 32'h0 : _GEN_865; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_867 = 10'h363 == _GEN_1280 ? 32'h0 : _GEN_866; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_868 = 10'h364 == _GEN_1280 ? 32'h0 : _GEN_867; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_869 = 10'h365 == _GEN_1280 ? 32'h0 : _GEN_868; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_870 = 10'h366 == _GEN_1280 ? 32'h0 : _GEN_869; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_871 = 10'h367 == _GEN_1280 ? 32'h0 : _GEN_870; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_872 = 10'h368 == _GEN_1280 ? 32'h0 : _GEN_871; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_873 = 10'h369 == _GEN_1280 ? 32'h0 : _GEN_872; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_874 = 10'h36a == _GEN_1280 ? 32'h0 : _GEN_873; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_875 = 10'h36b == _GEN_1280 ? 32'h0 : _GEN_874; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_876 = 10'h36c == _GEN_1280 ? 32'h0 : _GEN_875; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_877 = 10'h36d == _GEN_1280 ? 32'h0 : _GEN_876; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_878 = 10'h36e == _GEN_1280 ? 32'h0 : _GEN_877; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_879 = 10'h36f == _GEN_1280 ? 32'h0 : _GEN_878; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_880 = 10'h370 == _GEN_1280 ? 32'h0 : _GEN_879; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_881 = 10'h371 == _GEN_1280 ? 32'h0 : _GEN_880; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_882 = 10'h372 == _GEN_1280 ? 32'h0 : _GEN_881; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_883 = 10'h373 == _GEN_1280 ? 32'h0 : _GEN_882; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_884 = 10'h374 == _GEN_1280 ? 32'h0 : _GEN_883; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_885 = 10'h375 == _GEN_1280 ? 32'h0 : _GEN_884; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_886 = 10'h376 == _GEN_1280 ? 32'h0 : _GEN_885; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_887 = 10'h377 == _GEN_1280 ? 32'h0 : _GEN_886; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_888 = 10'h378 == _GEN_1280 ? 32'h0 : _GEN_887; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_889 = 10'h379 == _GEN_1280 ? 32'h0 : _GEN_888; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_890 = 10'h37a == _GEN_1280 ? 32'h0 : _GEN_889; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_891 = 10'h37b == _GEN_1280 ? 32'h0 : _GEN_890; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_892 = 10'h37c == _GEN_1280 ? 32'h0 : _GEN_891; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_893 = 10'h37d == _GEN_1280 ? 32'h0 : _GEN_892; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_894 = 10'h37e == _GEN_1280 ? 32'h0 : _GEN_893; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_895 = 10'h37f == _GEN_1280 ? 32'h0 : _GEN_894; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_896 = 10'h380 == _GEN_1280 ? 32'h0 : _GEN_895; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_897 = 10'h381 == _GEN_1280 ? 32'h0 : _GEN_896; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_898 = 10'h382 == _GEN_1280 ? 32'h0 : _GEN_897; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_899 = 10'h383 == _GEN_1280 ? 32'h0 : _GEN_898; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_900 = 10'h384 == _GEN_1280 ? 32'h0 : _GEN_899; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_901 = 10'h385 == _GEN_1280 ? 32'h0 : _GEN_900; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_902 = 10'h386 == _GEN_1280 ? 32'h0 : _GEN_901; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_903 = 10'h387 == _GEN_1280 ? 32'h0 : _GEN_902; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_904 = 10'h388 == _GEN_1280 ? 32'h0 : _GEN_903; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_905 = 10'h389 == _GEN_1280 ? 32'h0 : _GEN_904; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_906 = 10'h38a == _GEN_1280 ? 32'h0 : _GEN_905; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_907 = 10'h38b == _GEN_1280 ? 32'h0 : _GEN_906; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_908 = 10'h38c == _GEN_1280 ? 32'h0 : _GEN_907; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_909 = 10'h38d == _GEN_1280 ? 32'h0 : _GEN_908; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_910 = 10'h38e == _GEN_1280 ? 32'h0 : _GEN_909; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_911 = 10'h38f == _GEN_1280 ? 32'h0 : _GEN_910; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_912 = 10'h390 == _GEN_1280 ? 32'h0 : _GEN_911; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_913 = 10'h391 == _GEN_1280 ? 32'h0 : _GEN_912; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_914 = 10'h392 == _GEN_1280 ? 32'h0 : _GEN_913; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_915 = 10'h393 == _GEN_1280 ? 32'h0 : _GEN_914; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_916 = 10'h394 == _GEN_1280 ? 32'h0 : _GEN_915; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_917 = 10'h395 == _GEN_1280 ? 32'h0 : _GEN_916; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_918 = 10'h396 == _GEN_1280 ? 32'h0 : _GEN_917; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_919 = 10'h397 == _GEN_1280 ? 32'h0 : _GEN_918; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_920 = 10'h398 == _GEN_1280 ? 32'h0 : _GEN_919; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_921 = 10'h399 == _GEN_1280 ? 32'h0 : _GEN_920; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_922 = 10'h39a == _GEN_1280 ? 32'h0 : _GEN_921; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_923 = 10'h39b == _GEN_1280 ? 32'h0 : _GEN_922; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_924 = 10'h39c == _GEN_1280 ? 32'h0 : _GEN_923; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_925 = 10'h39d == _GEN_1280 ? 32'h0 : _GEN_924; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_926 = 10'h39e == _GEN_1280 ? 32'h0 : _GEN_925; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_927 = 10'h39f == _GEN_1280 ? 32'h0 : _GEN_926; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_928 = 10'h3a0 == _GEN_1280 ? 32'h0 : _GEN_927; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_929 = 10'h3a1 == _GEN_1280 ? 32'h0 : _GEN_928; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_930 = 10'h3a2 == _GEN_1280 ? 32'h0 : _GEN_929; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_931 = 10'h3a3 == _GEN_1280 ? 32'h0 : _GEN_930; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_932 = 10'h3a4 == _GEN_1280 ? 32'h0 : _GEN_931; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_933 = 10'h3a5 == _GEN_1280 ? 32'h0 : _GEN_932; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_934 = 10'h3a6 == _GEN_1280 ? 32'h0 : _GEN_933; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_935 = 10'h3a7 == _GEN_1280 ? 32'h0 : _GEN_934; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_936 = 10'h3a8 == _GEN_1280 ? 32'h0 : _GEN_935; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_937 = 10'h3a9 == _GEN_1280 ? 32'h0 : _GEN_936; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_938 = 10'h3aa == _GEN_1280 ? 32'h0 : _GEN_937; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_939 = 10'h3ab == _GEN_1280 ? 32'h0 : _GEN_938; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_940 = 10'h3ac == _GEN_1280 ? 32'h0 : _GEN_939; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_941 = 10'h3ad == _GEN_1280 ? 32'h0 : _GEN_940; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_942 = 10'h3ae == _GEN_1280 ? 32'h0 : _GEN_941; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_943 = 10'h3af == _GEN_1280 ? 32'h0 : _GEN_942; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_944 = 10'h3b0 == _GEN_1280 ? 32'h0 : _GEN_943; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_945 = 10'h3b1 == _GEN_1280 ? 32'h0 : _GEN_944; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_946 = 10'h3b2 == _GEN_1280 ? 32'h0 : _GEN_945; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_947 = 10'h3b3 == _GEN_1280 ? 32'h0 : _GEN_946; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_948 = 10'h3b4 == _GEN_1280 ? 32'h0 : _GEN_947; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_949 = 10'h3b5 == _GEN_1280 ? 32'h0 : _GEN_948; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_950 = 10'h3b6 == _GEN_1280 ? 32'h0 : _GEN_949; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_951 = 10'h3b7 == _GEN_1280 ? 32'h0 : _GEN_950; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_952 = 10'h3b8 == _GEN_1280 ? 32'h0 : _GEN_951; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_953 = 10'h3b9 == _GEN_1280 ? 32'h0 : _GEN_952; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_954 = 10'h3ba == _GEN_1280 ? 32'h0 : _GEN_953; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_955 = 10'h3bb == _GEN_1280 ? 32'h0 : _GEN_954; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_956 = 10'h3bc == _GEN_1280 ? 32'h0 : _GEN_955; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_957 = 10'h3bd == _GEN_1280 ? 32'h0 : _GEN_956; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_958 = 10'h3be == _GEN_1280 ? 32'h0 : _GEN_957; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_959 = 10'h3bf == _GEN_1280 ? 32'h0 : _GEN_958; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_960 = 10'h3c0 == _GEN_1280 ? 32'h0 : _GEN_959; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_961 = 10'h3c1 == _GEN_1280 ? 32'h0 : _GEN_960; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_962 = 10'h3c2 == _GEN_1280 ? 32'h0 : _GEN_961; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_963 = 10'h3c3 == _GEN_1280 ? 32'h0 : _GEN_962; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_964 = 10'h3c4 == _GEN_1280 ? 32'h0 : _GEN_963; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_965 = 10'h3c5 == _GEN_1280 ? 32'h0 : _GEN_964; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_966 = 10'h3c6 == _GEN_1280 ? 32'h0 : _GEN_965; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_967 = 10'h3c7 == _GEN_1280 ? 32'h0 : _GEN_966; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_968 = 10'h3c8 == _GEN_1280 ? 32'h0 : _GEN_967; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_969 = 10'h3c9 == _GEN_1280 ? 32'h0 : _GEN_968; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_970 = 10'h3ca == _GEN_1280 ? 32'h0 : _GEN_969; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_971 = 10'h3cb == _GEN_1280 ? 32'h0 : _GEN_970; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_972 = 10'h3cc == _GEN_1280 ? 32'h0 : _GEN_971; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_973 = 10'h3cd == _GEN_1280 ? 32'h0 : _GEN_972; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_974 = 10'h3ce == _GEN_1280 ? 32'h0 : _GEN_973; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_975 = 10'h3cf == _GEN_1280 ? 32'h0 : _GEN_974; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_976 = 10'h3d0 == _GEN_1280 ? 32'h0 : _GEN_975; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_977 = 10'h3d1 == _GEN_1280 ? 32'h0 : _GEN_976; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_978 = 10'h3d2 == _GEN_1280 ? 32'h0 : _GEN_977; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_979 = 10'h3d3 == _GEN_1280 ? 32'h0 : _GEN_978; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_980 = 10'h3d4 == _GEN_1280 ? 32'h0 : _GEN_979; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_981 = 10'h3d5 == _GEN_1280 ? 32'h0 : _GEN_980; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_982 = 10'h3d6 == _GEN_1280 ? 32'h0 : _GEN_981; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_983 = 10'h3d7 == _GEN_1280 ? 32'h0 : _GEN_982; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_984 = 10'h3d8 == _GEN_1280 ? 32'h0 : _GEN_983; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_985 = 10'h3d9 == _GEN_1280 ? 32'h0 : _GEN_984; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_986 = 10'h3da == _GEN_1280 ? 32'h0 : _GEN_985; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_987 = 10'h3db == _GEN_1280 ? 32'h0 : _GEN_986; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_988 = 10'h3dc == _GEN_1280 ? 32'h0 : _GEN_987; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_989 = 10'h3dd == _GEN_1280 ? 32'h0 : _GEN_988; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_990 = 10'h3de == _GEN_1280 ? 32'h0 : _GEN_989; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_991 = 10'h3df == _GEN_1280 ? 32'h0 : _GEN_990; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_992 = 10'h3e0 == _GEN_1280 ? 32'h0 : _GEN_991; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_993 = 10'h3e1 == _GEN_1280 ? 32'h0 : _GEN_992; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_994 = 10'h3e2 == _GEN_1280 ? 32'h0 : _GEN_993; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_995 = 10'h3e3 == _GEN_1280 ? 32'h0 : _GEN_994; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_996 = 10'h3e4 == _GEN_1280 ? 32'h0 : _GEN_995; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_997 = 10'h3e5 == _GEN_1280 ? 32'h0 : _GEN_996; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_998 = 10'h3e6 == _GEN_1280 ? 32'h0 : _GEN_997; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_999 = 10'h3e7 == _GEN_1280 ? 32'h0 : _GEN_998; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1000 = 10'h3e8 == _GEN_1280 ? 32'h0 : _GEN_999; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1001 = 10'h3e9 == _GEN_1280 ? 32'h0 : _GEN_1000; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1002 = 10'h3ea == _GEN_1280 ? 32'h0 : _GEN_1001; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1003 = 10'h3eb == _GEN_1280 ? 32'h0 : _GEN_1002; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1004 = 10'h3ec == _GEN_1280 ? 32'h0 : _GEN_1003; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1005 = 10'h3ed == _GEN_1280 ? 32'h0 : _GEN_1004; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1006 = 10'h3ee == _GEN_1280 ? 32'h0 : _GEN_1005; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1007 = 10'h3ef == _GEN_1280 ? 32'h0 : _GEN_1006; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1008 = 10'h3f0 == _GEN_1280 ? 32'h0 : _GEN_1007; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1009 = 10'h3f1 == _GEN_1280 ? 32'h0 : _GEN_1008; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1010 = 10'h3f2 == _GEN_1280 ? 32'h0 : _GEN_1009; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1011 = 10'h3f3 == _GEN_1280 ? 32'h0 : _GEN_1010; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1012 = 10'h3f4 == _GEN_1280 ? 32'h0 : _GEN_1011; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1013 = 10'h3f5 == _GEN_1280 ? 32'h0 : _GEN_1012; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1014 = 10'h3f6 == _GEN_1280 ? 32'h0 : _GEN_1013; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1015 = 10'h3f7 == _GEN_1280 ? 32'h0 : _GEN_1014; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1016 = 10'h3f8 == _GEN_1280 ? 32'h0 : _GEN_1015; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1017 = 10'h3f9 == _GEN_1280 ? 32'h0 : _GEN_1016; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1018 = 10'h3fa == _GEN_1280 ? 32'h0 : _GEN_1017; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1019 = 10'h3fb == _GEN_1280 ? 32'h0 : _GEN_1018; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1020 = 10'h3fc == _GEN_1280 ? 32'h0 : _GEN_1019; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1021 = 10'h3fd == _GEN_1280 ? 32'h0 : _GEN_1020; // @[InstMemory.scala 20:{11,11}]
  wire [31:0] _GEN_1022 = 10'h3fe == _GEN_1280 ? 32'h0 : _GEN_1021; // @[InstMemory.scala 20:{11,11}]
  assign io_inst = 10'h3ff == _GEN_1280 ? 32'h0 : _GEN_1022; // @[InstMemory.scala 20:{11,11}]
endmodule
module DData(
  input         clock,
  input         reset,
  input  [31:0] io_addr,
  input  [31:0] io_writeData,
  input         io_writeEnable,
  output [31:0] io_readData
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_0; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1; // @[DataMemory.scala 26:20]
  reg [31:0] ram_2; // @[DataMemory.scala 26:20]
  reg [31:0] ram_3; // @[DataMemory.scala 26:20]
  reg [31:0] ram_4; // @[DataMemory.scala 26:20]
  reg [31:0] ram_5; // @[DataMemory.scala 26:20]
  reg [31:0] ram_6; // @[DataMemory.scala 26:20]
  reg [31:0] ram_7; // @[DataMemory.scala 26:20]
  reg [31:0] ram_8; // @[DataMemory.scala 26:20]
  reg [31:0] ram_9; // @[DataMemory.scala 26:20]
  reg [31:0] ram_10; // @[DataMemory.scala 26:20]
  reg [31:0] ram_11; // @[DataMemory.scala 26:20]
  reg [31:0] ram_12; // @[DataMemory.scala 26:20]
  reg [31:0] ram_13; // @[DataMemory.scala 26:20]
  reg [31:0] ram_14; // @[DataMemory.scala 26:20]
  reg [31:0] ram_15; // @[DataMemory.scala 26:20]
  reg [31:0] ram_16; // @[DataMemory.scala 26:20]
  reg [31:0] ram_17; // @[DataMemory.scala 26:20]
  reg [31:0] ram_18; // @[DataMemory.scala 26:20]
  reg [31:0] ram_19; // @[DataMemory.scala 26:20]
  reg [31:0] ram_20; // @[DataMemory.scala 26:20]
  reg [31:0] ram_21; // @[DataMemory.scala 26:20]
  reg [31:0] ram_22; // @[DataMemory.scala 26:20]
  reg [31:0] ram_23; // @[DataMemory.scala 26:20]
  reg [31:0] ram_24; // @[DataMemory.scala 26:20]
  reg [31:0] ram_25; // @[DataMemory.scala 26:20]
  reg [31:0] ram_26; // @[DataMemory.scala 26:20]
  reg [31:0] ram_27; // @[DataMemory.scala 26:20]
  reg [31:0] ram_28; // @[DataMemory.scala 26:20]
  reg [31:0] ram_29; // @[DataMemory.scala 26:20]
  reg [31:0] ram_30; // @[DataMemory.scala 26:20]
  reg [31:0] ram_31; // @[DataMemory.scala 26:20]
  reg [31:0] ram_32; // @[DataMemory.scala 26:20]
  reg [31:0] ram_33; // @[DataMemory.scala 26:20]
  reg [31:0] ram_34; // @[DataMemory.scala 26:20]
  reg [31:0] ram_35; // @[DataMemory.scala 26:20]
  reg [31:0] ram_36; // @[DataMemory.scala 26:20]
  reg [31:0] ram_37; // @[DataMemory.scala 26:20]
  reg [31:0] ram_38; // @[DataMemory.scala 26:20]
  reg [31:0] ram_39; // @[DataMemory.scala 26:20]
  reg [31:0] ram_40; // @[DataMemory.scala 26:20]
  reg [31:0] ram_41; // @[DataMemory.scala 26:20]
  reg [31:0] ram_42; // @[DataMemory.scala 26:20]
  reg [31:0] ram_43; // @[DataMemory.scala 26:20]
  reg [31:0] ram_44; // @[DataMemory.scala 26:20]
  reg [31:0] ram_45; // @[DataMemory.scala 26:20]
  reg [31:0] ram_46; // @[DataMemory.scala 26:20]
  reg [31:0] ram_47; // @[DataMemory.scala 26:20]
  reg [31:0] ram_48; // @[DataMemory.scala 26:20]
  reg [31:0] ram_49; // @[DataMemory.scala 26:20]
  reg [31:0] ram_50; // @[DataMemory.scala 26:20]
  reg [31:0] ram_51; // @[DataMemory.scala 26:20]
  reg [31:0] ram_52; // @[DataMemory.scala 26:20]
  reg [31:0] ram_53; // @[DataMemory.scala 26:20]
  reg [31:0] ram_54; // @[DataMemory.scala 26:20]
  reg [31:0] ram_55; // @[DataMemory.scala 26:20]
  reg [31:0] ram_56; // @[DataMemory.scala 26:20]
  reg [31:0] ram_57; // @[DataMemory.scala 26:20]
  reg [31:0] ram_58; // @[DataMemory.scala 26:20]
  reg [31:0] ram_59; // @[DataMemory.scala 26:20]
  reg [31:0] ram_60; // @[DataMemory.scala 26:20]
  reg [31:0] ram_61; // @[DataMemory.scala 26:20]
  reg [31:0] ram_62; // @[DataMemory.scala 26:20]
  reg [31:0] ram_63; // @[DataMemory.scala 26:20]
  reg [31:0] ram_64; // @[DataMemory.scala 26:20]
  reg [31:0] ram_65; // @[DataMemory.scala 26:20]
  reg [31:0] ram_66; // @[DataMemory.scala 26:20]
  reg [31:0] ram_67; // @[DataMemory.scala 26:20]
  reg [31:0] ram_68; // @[DataMemory.scala 26:20]
  reg [31:0] ram_69; // @[DataMemory.scala 26:20]
  reg [31:0] ram_70; // @[DataMemory.scala 26:20]
  reg [31:0] ram_71; // @[DataMemory.scala 26:20]
  reg [31:0] ram_72; // @[DataMemory.scala 26:20]
  reg [31:0] ram_73; // @[DataMemory.scala 26:20]
  reg [31:0] ram_74; // @[DataMemory.scala 26:20]
  reg [31:0] ram_75; // @[DataMemory.scala 26:20]
  reg [31:0] ram_76; // @[DataMemory.scala 26:20]
  reg [31:0] ram_77; // @[DataMemory.scala 26:20]
  reg [31:0] ram_78; // @[DataMemory.scala 26:20]
  reg [31:0] ram_79; // @[DataMemory.scala 26:20]
  reg [31:0] ram_80; // @[DataMemory.scala 26:20]
  reg [31:0] ram_81; // @[DataMemory.scala 26:20]
  reg [31:0] ram_82; // @[DataMemory.scala 26:20]
  reg [31:0] ram_83; // @[DataMemory.scala 26:20]
  reg [31:0] ram_84; // @[DataMemory.scala 26:20]
  reg [31:0] ram_85; // @[DataMemory.scala 26:20]
  reg [31:0] ram_86; // @[DataMemory.scala 26:20]
  reg [31:0] ram_87; // @[DataMemory.scala 26:20]
  reg [31:0] ram_88; // @[DataMemory.scala 26:20]
  reg [31:0] ram_89; // @[DataMemory.scala 26:20]
  reg [31:0] ram_90; // @[DataMemory.scala 26:20]
  reg [31:0] ram_91; // @[DataMemory.scala 26:20]
  reg [31:0] ram_92; // @[DataMemory.scala 26:20]
  reg [31:0] ram_93; // @[DataMemory.scala 26:20]
  reg [31:0] ram_94; // @[DataMemory.scala 26:20]
  reg [31:0] ram_95; // @[DataMemory.scala 26:20]
  reg [31:0] ram_96; // @[DataMemory.scala 26:20]
  reg [31:0] ram_97; // @[DataMemory.scala 26:20]
  reg [31:0] ram_98; // @[DataMemory.scala 26:20]
  reg [31:0] ram_99; // @[DataMemory.scala 26:20]
  reg [31:0] ram_100; // @[DataMemory.scala 26:20]
  reg [31:0] ram_101; // @[DataMemory.scala 26:20]
  reg [31:0] ram_102; // @[DataMemory.scala 26:20]
  reg [31:0] ram_103; // @[DataMemory.scala 26:20]
  reg [31:0] ram_104; // @[DataMemory.scala 26:20]
  reg [31:0] ram_105; // @[DataMemory.scala 26:20]
  reg [31:0] ram_106; // @[DataMemory.scala 26:20]
  reg [31:0] ram_107; // @[DataMemory.scala 26:20]
  reg [31:0] ram_108; // @[DataMemory.scala 26:20]
  reg [31:0] ram_109; // @[DataMemory.scala 26:20]
  reg [31:0] ram_110; // @[DataMemory.scala 26:20]
  reg [31:0] ram_111; // @[DataMemory.scala 26:20]
  reg [31:0] ram_112; // @[DataMemory.scala 26:20]
  reg [31:0] ram_113; // @[DataMemory.scala 26:20]
  reg [31:0] ram_114; // @[DataMemory.scala 26:20]
  reg [31:0] ram_115; // @[DataMemory.scala 26:20]
  reg [31:0] ram_116; // @[DataMemory.scala 26:20]
  reg [31:0] ram_117; // @[DataMemory.scala 26:20]
  reg [31:0] ram_118; // @[DataMemory.scala 26:20]
  reg [31:0] ram_119; // @[DataMemory.scala 26:20]
  reg [31:0] ram_120; // @[DataMemory.scala 26:20]
  reg [31:0] ram_121; // @[DataMemory.scala 26:20]
  reg [31:0] ram_122; // @[DataMemory.scala 26:20]
  reg [31:0] ram_123; // @[DataMemory.scala 26:20]
  reg [31:0] ram_124; // @[DataMemory.scala 26:20]
  reg [31:0] ram_125; // @[DataMemory.scala 26:20]
  reg [31:0] ram_126; // @[DataMemory.scala 26:20]
  reg [31:0] ram_127; // @[DataMemory.scala 26:20]
  reg [31:0] ram_128; // @[DataMemory.scala 26:20]
  reg [31:0] ram_129; // @[DataMemory.scala 26:20]
  reg [31:0] ram_130; // @[DataMemory.scala 26:20]
  reg [31:0] ram_131; // @[DataMemory.scala 26:20]
  reg [31:0] ram_132; // @[DataMemory.scala 26:20]
  reg [31:0] ram_133; // @[DataMemory.scala 26:20]
  reg [31:0] ram_134; // @[DataMemory.scala 26:20]
  reg [31:0] ram_135; // @[DataMemory.scala 26:20]
  reg [31:0] ram_136; // @[DataMemory.scala 26:20]
  reg [31:0] ram_137; // @[DataMemory.scala 26:20]
  reg [31:0] ram_138; // @[DataMemory.scala 26:20]
  reg [31:0] ram_139; // @[DataMemory.scala 26:20]
  reg [31:0] ram_140; // @[DataMemory.scala 26:20]
  reg [31:0] ram_141; // @[DataMemory.scala 26:20]
  reg [31:0] ram_142; // @[DataMemory.scala 26:20]
  reg [31:0] ram_143; // @[DataMemory.scala 26:20]
  reg [31:0] ram_144; // @[DataMemory.scala 26:20]
  reg [31:0] ram_145; // @[DataMemory.scala 26:20]
  reg [31:0] ram_146; // @[DataMemory.scala 26:20]
  reg [31:0] ram_147; // @[DataMemory.scala 26:20]
  reg [31:0] ram_148; // @[DataMemory.scala 26:20]
  reg [31:0] ram_149; // @[DataMemory.scala 26:20]
  reg [31:0] ram_150; // @[DataMemory.scala 26:20]
  reg [31:0] ram_151; // @[DataMemory.scala 26:20]
  reg [31:0] ram_152; // @[DataMemory.scala 26:20]
  reg [31:0] ram_153; // @[DataMemory.scala 26:20]
  reg [31:0] ram_154; // @[DataMemory.scala 26:20]
  reg [31:0] ram_155; // @[DataMemory.scala 26:20]
  reg [31:0] ram_156; // @[DataMemory.scala 26:20]
  reg [31:0] ram_157; // @[DataMemory.scala 26:20]
  reg [31:0] ram_158; // @[DataMemory.scala 26:20]
  reg [31:0] ram_159; // @[DataMemory.scala 26:20]
  reg [31:0] ram_160; // @[DataMemory.scala 26:20]
  reg [31:0] ram_161; // @[DataMemory.scala 26:20]
  reg [31:0] ram_162; // @[DataMemory.scala 26:20]
  reg [31:0] ram_163; // @[DataMemory.scala 26:20]
  reg [31:0] ram_164; // @[DataMemory.scala 26:20]
  reg [31:0] ram_165; // @[DataMemory.scala 26:20]
  reg [31:0] ram_166; // @[DataMemory.scala 26:20]
  reg [31:0] ram_167; // @[DataMemory.scala 26:20]
  reg [31:0] ram_168; // @[DataMemory.scala 26:20]
  reg [31:0] ram_169; // @[DataMemory.scala 26:20]
  reg [31:0] ram_170; // @[DataMemory.scala 26:20]
  reg [31:0] ram_171; // @[DataMemory.scala 26:20]
  reg [31:0] ram_172; // @[DataMemory.scala 26:20]
  reg [31:0] ram_173; // @[DataMemory.scala 26:20]
  reg [31:0] ram_174; // @[DataMemory.scala 26:20]
  reg [31:0] ram_175; // @[DataMemory.scala 26:20]
  reg [31:0] ram_176; // @[DataMemory.scala 26:20]
  reg [31:0] ram_177; // @[DataMemory.scala 26:20]
  reg [31:0] ram_178; // @[DataMemory.scala 26:20]
  reg [31:0] ram_179; // @[DataMemory.scala 26:20]
  reg [31:0] ram_180; // @[DataMemory.scala 26:20]
  reg [31:0] ram_181; // @[DataMemory.scala 26:20]
  reg [31:0] ram_182; // @[DataMemory.scala 26:20]
  reg [31:0] ram_183; // @[DataMemory.scala 26:20]
  reg [31:0] ram_184; // @[DataMemory.scala 26:20]
  reg [31:0] ram_185; // @[DataMemory.scala 26:20]
  reg [31:0] ram_186; // @[DataMemory.scala 26:20]
  reg [31:0] ram_187; // @[DataMemory.scala 26:20]
  reg [31:0] ram_188; // @[DataMemory.scala 26:20]
  reg [31:0] ram_189; // @[DataMemory.scala 26:20]
  reg [31:0] ram_190; // @[DataMemory.scala 26:20]
  reg [31:0] ram_191; // @[DataMemory.scala 26:20]
  reg [31:0] ram_192; // @[DataMemory.scala 26:20]
  reg [31:0] ram_193; // @[DataMemory.scala 26:20]
  reg [31:0] ram_194; // @[DataMemory.scala 26:20]
  reg [31:0] ram_195; // @[DataMemory.scala 26:20]
  reg [31:0] ram_196; // @[DataMemory.scala 26:20]
  reg [31:0] ram_197; // @[DataMemory.scala 26:20]
  reg [31:0] ram_198; // @[DataMemory.scala 26:20]
  reg [31:0] ram_199; // @[DataMemory.scala 26:20]
  reg [31:0] ram_200; // @[DataMemory.scala 26:20]
  reg [31:0] ram_201; // @[DataMemory.scala 26:20]
  reg [31:0] ram_202; // @[DataMemory.scala 26:20]
  reg [31:0] ram_203; // @[DataMemory.scala 26:20]
  reg [31:0] ram_204; // @[DataMemory.scala 26:20]
  reg [31:0] ram_205; // @[DataMemory.scala 26:20]
  reg [31:0] ram_206; // @[DataMemory.scala 26:20]
  reg [31:0] ram_207; // @[DataMemory.scala 26:20]
  reg [31:0] ram_208; // @[DataMemory.scala 26:20]
  reg [31:0] ram_209; // @[DataMemory.scala 26:20]
  reg [31:0] ram_210; // @[DataMemory.scala 26:20]
  reg [31:0] ram_211; // @[DataMemory.scala 26:20]
  reg [31:0] ram_212; // @[DataMemory.scala 26:20]
  reg [31:0] ram_213; // @[DataMemory.scala 26:20]
  reg [31:0] ram_214; // @[DataMemory.scala 26:20]
  reg [31:0] ram_215; // @[DataMemory.scala 26:20]
  reg [31:0] ram_216; // @[DataMemory.scala 26:20]
  reg [31:0] ram_217; // @[DataMemory.scala 26:20]
  reg [31:0] ram_218; // @[DataMemory.scala 26:20]
  reg [31:0] ram_219; // @[DataMemory.scala 26:20]
  reg [31:0] ram_220; // @[DataMemory.scala 26:20]
  reg [31:0] ram_221; // @[DataMemory.scala 26:20]
  reg [31:0] ram_222; // @[DataMemory.scala 26:20]
  reg [31:0] ram_223; // @[DataMemory.scala 26:20]
  reg [31:0] ram_224; // @[DataMemory.scala 26:20]
  reg [31:0] ram_225; // @[DataMemory.scala 26:20]
  reg [31:0] ram_226; // @[DataMemory.scala 26:20]
  reg [31:0] ram_227; // @[DataMemory.scala 26:20]
  reg [31:0] ram_228; // @[DataMemory.scala 26:20]
  reg [31:0] ram_229; // @[DataMemory.scala 26:20]
  reg [31:0] ram_230; // @[DataMemory.scala 26:20]
  reg [31:0] ram_231; // @[DataMemory.scala 26:20]
  reg [31:0] ram_232; // @[DataMemory.scala 26:20]
  reg [31:0] ram_233; // @[DataMemory.scala 26:20]
  reg [31:0] ram_234; // @[DataMemory.scala 26:20]
  reg [31:0] ram_235; // @[DataMemory.scala 26:20]
  reg [31:0] ram_236; // @[DataMemory.scala 26:20]
  reg [31:0] ram_237; // @[DataMemory.scala 26:20]
  reg [31:0] ram_238; // @[DataMemory.scala 26:20]
  reg [31:0] ram_239; // @[DataMemory.scala 26:20]
  reg [31:0] ram_240; // @[DataMemory.scala 26:20]
  reg [31:0] ram_241; // @[DataMemory.scala 26:20]
  reg [31:0] ram_242; // @[DataMemory.scala 26:20]
  reg [31:0] ram_243; // @[DataMemory.scala 26:20]
  reg [31:0] ram_244; // @[DataMemory.scala 26:20]
  reg [31:0] ram_245; // @[DataMemory.scala 26:20]
  reg [31:0] ram_246; // @[DataMemory.scala 26:20]
  reg [31:0] ram_247; // @[DataMemory.scala 26:20]
  reg [31:0] ram_248; // @[DataMemory.scala 26:20]
  reg [31:0] ram_249; // @[DataMemory.scala 26:20]
  reg [31:0] ram_250; // @[DataMemory.scala 26:20]
  reg [31:0] ram_251; // @[DataMemory.scala 26:20]
  reg [31:0] ram_252; // @[DataMemory.scala 26:20]
  reg [31:0] ram_253; // @[DataMemory.scala 26:20]
  reg [31:0] ram_254; // @[DataMemory.scala 26:20]
  reg [31:0] ram_255; // @[DataMemory.scala 26:20]
  reg [31:0] ram_256; // @[DataMemory.scala 26:20]
  reg [31:0] ram_257; // @[DataMemory.scala 26:20]
  reg [31:0] ram_258; // @[DataMemory.scala 26:20]
  reg [31:0] ram_259; // @[DataMemory.scala 26:20]
  reg [31:0] ram_260; // @[DataMemory.scala 26:20]
  reg [31:0] ram_261; // @[DataMemory.scala 26:20]
  reg [31:0] ram_262; // @[DataMemory.scala 26:20]
  reg [31:0] ram_263; // @[DataMemory.scala 26:20]
  reg [31:0] ram_264; // @[DataMemory.scala 26:20]
  reg [31:0] ram_265; // @[DataMemory.scala 26:20]
  reg [31:0] ram_266; // @[DataMemory.scala 26:20]
  reg [31:0] ram_267; // @[DataMemory.scala 26:20]
  reg [31:0] ram_268; // @[DataMemory.scala 26:20]
  reg [31:0] ram_269; // @[DataMemory.scala 26:20]
  reg [31:0] ram_270; // @[DataMemory.scala 26:20]
  reg [31:0] ram_271; // @[DataMemory.scala 26:20]
  reg [31:0] ram_272; // @[DataMemory.scala 26:20]
  reg [31:0] ram_273; // @[DataMemory.scala 26:20]
  reg [31:0] ram_274; // @[DataMemory.scala 26:20]
  reg [31:0] ram_275; // @[DataMemory.scala 26:20]
  reg [31:0] ram_276; // @[DataMemory.scala 26:20]
  reg [31:0] ram_277; // @[DataMemory.scala 26:20]
  reg [31:0] ram_278; // @[DataMemory.scala 26:20]
  reg [31:0] ram_279; // @[DataMemory.scala 26:20]
  reg [31:0] ram_280; // @[DataMemory.scala 26:20]
  reg [31:0] ram_281; // @[DataMemory.scala 26:20]
  reg [31:0] ram_282; // @[DataMemory.scala 26:20]
  reg [31:0] ram_283; // @[DataMemory.scala 26:20]
  reg [31:0] ram_284; // @[DataMemory.scala 26:20]
  reg [31:0] ram_285; // @[DataMemory.scala 26:20]
  reg [31:0] ram_286; // @[DataMemory.scala 26:20]
  reg [31:0] ram_287; // @[DataMemory.scala 26:20]
  reg [31:0] ram_288; // @[DataMemory.scala 26:20]
  reg [31:0] ram_289; // @[DataMemory.scala 26:20]
  reg [31:0] ram_290; // @[DataMemory.scala 26:20]
  reg [31:0] ram_291; // @[DataMemory.scala 26:20]
  reg [31:0] ram_292; // @[DataMemory.scala 26:20]
  reg [31:0] ram_293; // @[DataMemory.scala 26:20]
  reg [31:0] ram_294; // @[DataMemory.scala 26:20]
  reg [31:0] ram_295; // @[DataMemory.scala 26:20]
  reg [31:0] ram_296; // @[DataMemory.scala 26:20]
  reg [31:0] ram_297; // @[DataMemory.scala 26:20]
  reg [31:0] ram_298; // @[DataMemory.scala 26:20]
  reg [31:0] ram_299; // @[DataMemory.scala 26:20]
  reg [31:0] ram_300; // @[DataMemory.scala 26:20]
  reg [31:0] ram_301; // @[DataMemory.scala 26:20]
  reg [31:0] ram_302; // @[DataMemory.scala 26:20]
  reg [31:0] ram_303; // @[DataMemory.scala 26:20]
  reg [31:0] ram_304; // @[DataMemory.scala 26:20]
  reg [31:0] ram_305; // @[DataMemory.scala 26:20]
  reg [31:0] ram_306; // @[DataMemory.scala 26:20]
  reg [31:0] ram_307; // @[DataMemory.scala 26:20]
  reg [31:0] ram_308; // @[DataMemory.scala 26:20]
  reg [31:0] ram_309; // @[DataMemory.scala 26:20]
  reg [31:0] ram_310; // @[DataMemory.scala 26:20]
  reg [31:0] ram_311; // @[DataMemory.scala 26:20]
  reg [31:0] ram_312; // @[DataMemory.scala 26:20]
  reg [31:0] ram_313; // @[DataMemory.scala 26:20]
  reg [31:0] ram_314; // @[DataMemory.scala 26:20]
  reg [31:0] ram_315; // @[DataMemory.scala 26:20]
  reg [31:0] ram_316; // @[DataMemory.scala 26:20]
  reg [31:0] ram_317; // @[DataMemory.scala 26:20]
  reg [31:0] ram_318; // @[DataMemory.scala 26:20]
  reg [31:0] ram_319; // @[DataMemory.scala 26:20]
  reg [31:0] ram_320; // @[DataMemory.scala 26:20]
  reg [31:0] ram_321; // @[DataMemory.scala 26:20]
  reg [31:0] ram_322; // @[DataMemory.scala 26:20]
  reg [31:0] ram_323; // @[DataMemory.scala 26:20]
  reg [31:0] ram_324; // @[DataMemory.scala 26:20]
  reg [31:0] ram_325; // @[DataMemory.scala 26:20]
  reg [31:0] ram_326; // @[DataMemory.scala 26:20]
  reg [31:0] ram_327; // @[DataMemory.scala 26:20]
  reg [31:0] ram_328; // @[DataMemory.scala 26:20]
  reg [31:0] ram_329; // @[DataMemory.scala 26:20]
  reg [31:0] ram_330; // @[DataMemory.scala 26:20]
  reg [31:0] ram_331; // @[DataMemory.scala 26:20]
  reg [31:0] ram_332; // @[DataMemory.scala 26:20]
  reg [31:0] ram_333; // @[DataMemory.scala 26:20]
  reg [31:0] ram_334; // @[DataMemory.scala 26:20]
  reg [31:0] ram_335; // @[DataMemory.scala 26:20]
  reg [31:0] ram_336; // @[DataMemory.scala 26:20]
  reg [31:0] ram_337; // @[DataMemory.scala 26:20]
  reg [31:0] ram_338; // @[DataMemory.scala 26:20]
  reg [31:0] ram_339; // @[DataMemory.scala 26:20]
  reg [31:0] ram_340; // @[DataMemory.scala 26:20]
  reg [31:0] ram_341; // @[DataMemory.scala 26:20]
  reg [31:0] ram_342; // @[DataMemory.scala 26:20]
  reg [31:0] ram_343; // @[DataMemory.scala 26:20]
  reg [31:0] ram_344; // @[DataMemory.scala 26:20]
  reg [31:0] ram_345; // @[DataMemory.scala 26:20]
  reg [31:0] ram_346; // @[DataMemory.scala 26:20]
  reg [31:0] ram_347; // @[DataMemory.scala 26:20]
  reg [31:0] ram_348; // @[DataMemory.scala 26:20]
  reg [31:0] ram_349; // @[DataMemory.scala 26:20]
  reg [31:0] ram_350; // @[DataMemory.scala 26:20]
  reg [31:0] ram_351; // @[DataMemory.scala 26:20]
  reg [31:0] ram_352; // @[DataMemory.scala 26:20]
  reg [31:0] ram_353; // @[DataMemory.scala 26:20]
  reg [31:0] ram_354; // @[DataMemory.scala 26:20]
  reg [31:0] ram_355; // @[DataMemory.scala 26:20]
  reg [31:0] ram_356; // @[DataMemory.scala 26:20]
  reg [31:0] ram_357; // @[DataMemory.scala 26:20]
  reg [31:0] ram_358; // @[DataMemory.scala 26:20]
  reg [31:0] ram_359; // @[DataMemory.scala 26:20]
  reg [31:0] ram_360; // @[DataMemory.scala 26:20]
  reg [31:0] ram_361; // @[DataMemory.scala 26:20]
  reg [31:0] ram_362; // @[DataMemory.scala 26:20]
  reg [31:0] ram_363; // @[DataMemory.scala 26:20]
  reg [31:0] ram_364; // @[DataMemory.scala 26:20]
  reg [31:0] ram_365; // @[DataMemory.scala 26:20]
  reg [31:0] ram_366; // @[DataMemory.scala 26:20]
  reg [31:0] ram_367; // @[DataMemory.scala 26:20]
  reg [31:0] ram_368; // @[DataMemory.scala 26:20]
  reg [31:0] ram_369; // @[DataMemory.scala 26:20]
  reg [31:0] ram_370; // @[DataMemory.scala 26:20]
  reg [31:0] ram_371; // @[DataMemory.scala 26:20]
  reg [31:0] ram_372; // @[DataMemory.scala 26:20]
  reg [31:0] ram_373; // @[DataMemory.scala 26:20]
  reg [31:0] ram_374; // @[DataMemory.scala 26:20]
  reg [31:0] ram_375; // @[DataMemory.scala 26:20]
  reg [31:0] ram_376; // @[DataMemory.scala 26:20]
  reg [31:0] ram_377; // @[DataMemory.scala 26:20]
  reg [31:0] ram_378; // @[DataMemory.scala 26:20]
  reg [31:0] ram_379; // @[DataMemory.scala 26:20]
  reg [31:0] ram_380; // @[DataMemory.scala 26:20]
  reg [31:0] ram_381; // @[DataMemory.scala 26:20]
  reg [31:0] ram_382; // @[DataMemory.scala 26:20]
  reg [31:0] ram_383; // @[DataMemory.scala 26:20]
  reg [31:0] ram_384; // @[DataMemory.scala 26:20]
  reg [31:0] ram_385; // @[DataMemory.scala 26:20]
  reg [31:0] ram_386; // @[DataMemory.scala 26:20]
  reg [31:0] ram_387; // @[DataMemory.scala 26:20]
  reg [31:0] ram_388; // @[DataMemory.scala 26:20]
  reg [31:0] ram_389; // @[DataMemory.scala 26:20]
  reg [31:0] ram_390; // @[DataMemory.scala 26:20]
  reg [31:0] ram_391; // @[DataMemory.scala 26:20]
  reg [31:0] ram_392; // @[DataMemory.scala 26:20]
  reg [31:0] ram_393; // @[DataMemory.scala 26:20]
  reg [31:0] ram_394; // @[DataMemory.scala 26:20]
  reg [31:0] ram_395; // @[DataMemory.scala 26:20]
  reg [31:0] ram_396; // @[DataMemory.scala 26:20]
  reg [31:0] ram_397; // @[DataMemory.scala 26:20]
  reg [31:0] ram_398; // @[DataMemory.scala 26:20]
  reg [31:0] ram_399; // @[DataMemory.scala 26:20]
  reg [31:0] ram_400; // @[DataMemory.scala 26:20]
  reg [31:0] ram_401; // @[DataMemory.scala 26:20]
  reg [31:0] ram_402; // @[DataMemory.scala 26:20]
  reg [31:0] ram_403; // @[DataMemory.scala 26:20]
  reg [31:0] ram_404; // @[DataMemory.scala 26:20]
  reg [31:0] ram_405; // @[DataMemory.scala 26:20]
  reg [31:0] ram_406; // @[DataMemory.scala 26:20]
  reg [31:0] ram_407; // @[DataMemory.scala 26:20]
  reg [31:0] ram_408; // @[DataMemory.scala 26:20]
  reg [31:0] ram_409; // @[DataMemory.scala 26:20]
  reg [31:0] ram_410; // @[DataMemory.scala 26:20]
  reg [31:0] ram_411; // @[DataMemory.scala 26:20]
  reg [31:0] ram_412; // @[DataMemory.scala 26:20]
  reg [31:0] ram_413; // @[DataMemory.scala 26:20]
  reg [31:0] ram_414; // @[DataMemory.scala 26:20]
  reg [31:0] ram_415; // @[DataMemory.scala 26:20]
  reg [31:0] ram_416; // @[DataMemory.scala 26:20]
  reg [31:0] ram_417; // @[DataMemory.scala 26:20]
  reg [31:0] ram_418; // @[DataMemory.scala 26:20]
  reg [31:0] ram_419; // @[DataMemory.scala 26:20]
  reg [31:0] ram_420; // @[DataMemory.scala 26:20]
  reg [31:0] ram_421; // @[DataMemory.scala 26:20]
  reg [31:0] ram_422; // @[DataMemory.scala 26:20]
  reg [31:0] ram_423; // @[DataMemory.scala 26:20]
  reg [31:0] ram_424; // @[DataMemory.scala 26:20]
  reg [31:0] ram_425; // @[DataMemory.scala 26:20]
  reg [31:0] ram_426; // @[DataMemory.scala 26:20]
  reg [31:0] ram_427; // @[DataMemory.scala 26:20]
  reg [31:0] ram_428; // @[DataMemory.scala 26:20]
  reg [31:0] ram_429; // @[DataMemory.scala 26:20]
  reg [31:0] ram_430; // @[DataMemory.scala 26:20]
  reg [31:0] ram_431; // @[DataMemory.scala 26:20]
  reg [31:0] ram_432; // @[DataMemory.scala 26:20]
  reg [31:0] ram_433; // @[DataMemory.scala 26:20]
  reg [31:0] ram_434; // @[DataMemory.scala 26:20]
  reg [31:0] ram_435; // @[DataMemory.scala 26:20]
  reg [31:0] ram_436; // @[DataMemory.scala 26:20]
  reg [31:0] ram_437; // @[DataMemory.scala 26:20]
  reg [31:0] ram_438; // @[DataMemory.scala 26:20]
  reg [31:0] ram_439; // @[DataMemory.scala 26:20]
  reg [31:0] ram_440; // @[DataMemory.scala 26:20]
  reg [31:0] ram_441; // @[DataMemory.scala 26:20]
  reg [31:0] ram_442; // @[DataMemory.scala 26:20]
  reg [31:0] ram_443; // @[DataMemory.scala 26:20]
  reg [31:0] ram_444; // @[DataMemory.scala 26:20]
  reg [31:0] ram_445; // @[DataMemory.scala 26:20]
  reg [31:0] ram_446; // @[DataMemory.scala 26:20]
  reg [31:0] ram_447; // @[DataMemory.scala 26:20]
  reg [31:0] ram_448; // @[DataMemory.scala 26:20]
  reg [31:0] ram_449; // @[DataMemory.scala 26:20]
  reg [31:0] ram_450; // @[DataMemory.scala 26:20]
  reg [31:0] ram_451; // @[DataMemory.scala 26:20]
  reg [31:0] ram_452; // @[DataMemory.scala 26:20]
  reg [31:0] ram_453; // @[DataMemory.scala 26:20]
  reg [31:0] ram_454; // @[DataMemory.scala 26:20]
  reg [31:0] ram_455; // @[DataMemory.scala 26:20]
  reg [31:0] ram_456; // @[DataMemory.scala 26:20]
  reg [31:0] ram_457; // @[DataMemory.scala 26:20]
  reg [31:0] ram_458; // @[DataMemory.scala 26:20]
  reg [31:0] ram_459; // @[DataMemory.scala 26:20]
  reg [31:0] ram_460; // @[DataMemory.scala 26:20]
  reg [31:0] ram_461; // @[DataMemory.scala 26:20]
  reg [31:0] ram_462; // @[DataMemory.scala 26:20]
  reg [31:0] ram_463; // @[DataMemory.scala 26:20]
  reg [31:0] ram_464; // @[DataMemory.scala 26:20]
  reg [31:0] ram_465; // @[DataMemory.scala 26:20]
  reg [31:0] ram_466; // @[DataMemory.scala 26:20]
  reg [31:0] ram_467; // @[DataMemory.scala 26:20]
  reg [31:0] ram_468; // @[DataMemory.scala 26:20]
  reg [31:0] ram_469; // @[DataMemory.scala 26:20]
  reg [31:0] ram_470; // @[DataMemory.scala 26:20]
  reg [31:0] ram_471; // @[DataMemory.scala 26:20]
  reg [31:0] ram_472; // @[DataMemory.scala 26:20]
  reg [31:0] ram_473; // @[DataMemory.scala 26:20]
  reg [31:0] ram_474; // @[DataMemory.scala 26:20]
  reg [31:0] ram_475; // @[DataMemory.scala 26:20]
  reg [31:0] ram_476; // @[DataMemory.scala 26:20]
  reg [31:0] ram_477; // @[DataMemory.scala 26:20]
  reg [31:0] ram_478; // @[DataMemory.scala 26:20]
  reg [31:0] ram_479; // @[DataMemory.scala 26:20]
  reg [31:0] ram_480; // @[DataMemory.scala 26:20]
  reg [31:0] ram_481; // @[DataMemory.scala 26:20]
  reg [31:0] ram_482; // @[DataMemory.scala 26:20]
  reg [31:0] ram_483; // @[DataMemory.scala 26:20]
  reg [31:0] ram_484; // @[DataMemory.scala 26:20]
  reg [31:0] ram_485; // @[DataMemory.scala 26:20]
  reg [31:0] ram_486; // @[DataMemory.scala 26:20]
  reg [31:0] ram_487; // @[DataMemory.scala 26:20]
  reg [31:0] ram_488; // @[DataMemory.scala 26:20]
  reg [31:0] ram_489; // @[DataMemory.scala 26:20]
  reg [31:0] ram_490; // @[DataMemory.scala 26:20]
  reg [31:0] ram_491; // @[DataMemory.scala 26:20]
  reg [31:0] ram_492; // @[DataMemory.scala 26:20]
  reg [31:0] ram_493; // @[DataMemory.scala 26:20]
  reg [31:0] ram_494; // @[DataMemory.scala 26:20]
  reg [31:0] ram_495; // @[DataMemory.scala 26:20]
  reg [31:0] ram_496; // @[DataMemory.scala 26:20]
  reg [31:0] ram_497; // @[DataMemory.scala 26:20]
  reg [31:0] ram_498; // @[DataMemory.scala 26:20]
  reg [31:0] ram_499; // @[DataMemory.scala 26:20]
  reg [31:0] ram_500; // @[DataMemory.scala 26:20]
  reg [31:0] ram_501; // @[DataMemory.scala 26:20]
  reg [31:0] ram_502; // @[DataMemory.scala 26:20]
  reg [31:0] ram_503; // @[DataMemory.scala 26:20]
  reg [31:0] ram_504; // @[DataMemory.scala 26:20]
  reg [31:0] ram_505; // @[DataMemory.scala 26:20]
  reg [31:0] ram_506; // @[DataMemory.scala 26:20]
  reg [31:0] ram_507; // @[DataMemory.scala 26:20]
  reg [31:0] ram_508; // @[DataMemory.scala 26:20]
  reg [31:0] ram_509; // @[DataMemory.scala 26:20]
  reg [31:0] ram_510; // @[DataMemory.scala 26:20]
  reg [31:0] ram_511; // @[DataMemory.scala 26:20]
  reg [31:0] ram_512; // @[DataMemory.scala 26:20]
  reg [31:0] ram_513; // @[DataMemory.scala 26:20]
  reg [31:0] ram_514; // @[DataMemory.scala 26:20]
  reg [31:0] ram_515; // @[DataMemory.scala 26:20]
  reg [31:0] ram_516; // @[DataMemory.scala 26:20]
  reg [31:0] ram_517; // @[DataMemory.scala 26:20]
  reg [31:0] ram_518; // @[DataMemory.scala 26:20]
  reg [31:0] ram_519; // @[DataMemory.scala 26:20]
  reg [31:0] ram_520; // @[DataMemory.scala 26:20]
  reg [31:0] ram_521; // @[DataMemory.scala 26:20]
  reg [31:0] ram_522; // @[DataMemory.scala 26:20]
  reg [31:0] ram_523; // @[DataMemory.scala 26:20]
  reg [31:0] ram_524; // @[DataMemory.scala 26:20]
  reg [31:0] ram_525; // @[DataMemory.scala 26:20]
  reg [31:0] ram_526; // @[DataMemory.scala 26:20]
  reg [31:0] ram_527; // @[DataMemory.scala 26:20]
  reg [31:0] ram_528; // @[DataMemory.scala 26:20]
  reg [31:0] ram_529; // @[DataMemory.scala 26:20]
  reg [31:0] ram_530; // @[DataMemory.scala 26:20]
  reg [31:0] ram_531; // @[DataMemory.scala 26:20]
  reg [31:0] ram_532; // @[DataMemory.scala 26:20]
  reg [31:0] ram_533; // @[DataMemory.scala 26:20]
  reg [31:0] ram_534; // @[DataMemory.scala 26:20]
  reg [31:0] ram_535; // @[DataMemory.scala 26:20]
  reg [31:0] ram_536; // @[DataMemory.scala 26:20]
  reg [31:0] ram_537; // @[DataMemory.scala 26:20]
  reg [31:0] ram_538; // @[DataMemory.scala 26:20]
  reg [31:0] ram_539; // @[DataMemory.scala 26:20]
  reg [31:0] ram_540; // @[DataMemory.scala 26:20]
  reg [31:0] ram_541; // @[DataMemory.scala 26:20]
  reg [31:0] ram_542; // @[DataMemory.scala 26:20]
  reg [31:0] ram_543; // @[DataMemory.scala 26:20]
  reg [31:0] ram_544; // @[DataMemory.scala 26:20]
  reg [31:0] ram_545; // @[DataMemory.scala 26:20]
  reg [31:0] ram_546; // @[DataMemory.scala 26:20]
  reg [31:0] ram_547; // @[DataMemory.scala 26:20]
  reg [31:0] ram_548; // @[DataMemory.scala 26:20]
  reg [31:0] ram_549; // @[DataMemory.scala 26:20]
  reg [31:0] ram_550; // @[DataMemory.scala 26:20]
  reg [31:0] ram_551; // @[DataMemory.scala 26:20]
  reg [31:0] ram_552; // @[DataMemory.scala 26:20]
  reg [31:0] ram_553; // @[DataMemory.scala 26:20]
  reg [31:0] ram_554; // @[DataMemory.scala 26:20]
  reg [31:0] ram_555; // @[DataMemory.scala 26:20]
  reg [31:0] ram_556; // @[DataMemory.scala 26:20]
  reg [31:0] ram_557; // @[DataMemory.scala 26:20]
  reg [31:0] ram_558; // @[DataMemory.scala 26:20]
  reg [31:0] ram_559; // @[DataMemory.scala 26:20]
  reg [31:0] ram_560; // @[DataMemory.scala 26:20]
  reg [31:0] ram_561; // @[DataMemory.scala 26:20]
  reg [31:0] ram_562; // @[DataMemory.scala 26:20]
  reg [31:0] ram_563; // @[DataMemory.scala 26:20]
  reg [31:0] ram_564; // @[DataMemory.scala 26:20]
  reg [31:0] ram_565; // @[DataMemory.scala 26:20]
  reg [31:0] ram_566; // @[DataMemory.scala 26:20]
  reg [31:0] ram_567; // @[DataMemory.scala 26:20]
  reg [31:0] ram_568; // @[DataMemory.scala 26:20]
  reg [31:0] ram_569; // @[DataMemory.scala 26:20]
  reg [31:0] ram_570; // @[DataMemory.scala 26:20]
  reg [31:0] ram_571; // @[DataMemory.scala 26:20]
  reg [31:0] ram_572; // @[DataMemory.scala 26:20]
  reg [31:0] ram_573; // @[DataMemory.scala 26:20]
  reg [31:0] ram_574; // @[DataMemory.scala 26:20]
  reg [31:0] ram_575; // @[DataMemory.scala 26:20]
  reg [31:0] ram_576; // @[DataMemory.scala 26:20]
  reg [31:0] ram_577; // @[DataMemory.scala 26:20]
  reg [31:0] ram_578; // @[DataMemory.scala 26:20]
  reg [31:0] ram_579; // @[DataMemory.scala 26:20]
  reg [31:0] ram_580; // @[DataMemory.scala 26:20]
  reg [31:0] ram_581; // @[DataMemory.scala 26:20]
  reg [31:0] ram_582; // @[DataMemory.scala 26:20]
  reg [31:0] ram_583; // @[DataMemory.scala 26:20]
  reg [31:0] ram_584; // @[DataMemory.scala 26:20]
  reg [31:0] ram_585; // @[DataMemory.scala 26:20]
  reg [31:0] ram_586; // @[DataMemory.scala 26:20]
  reg [31:0] ram_587; // @[DataMemory.scala 26:20]
  reg [31:0] ram_588; // @[DataMemory.scala 26:20]
  reg [31:0] ram_589; // @[DataMemory.scala 26:20]
  reg [31:0] ram_590; // @[DataMemory.scala 26:20]
  reg [31:0] ram_591; // @[DataMemory.scala 26:20]
  reg [31:0] ram_592; // @[DataMemory.scala 26:20]
  reg [31:0] ram_593; // @[DataMemory.scala 26:20]
  reg [31:0] ram_594; // @[DataMemory.scala 26:20]
  reg [31:0] ram_595; // @[DataMemory.scala 26:20]
  reg [31:0] ram_596; // @[DataMemory.scala 26:20]
  reg [31:0] ram_597; // @[DataMemory.scala 26:20]
  reg [31:0] ram_598; // @[DataMemory.scala 26:20]
  reg [31:0] ram_599; // @[DataMemory.scala 26:20]
  reg [31:0] ram_600; // @[DataMemory.scala 26:20]
  reg [31:0] ram_601; // @[DataMemory.scala 26:20]
  reg [31:0] ram_602; // @[DataMemory.scala 26:20]
  reg [31:0] ram_603; // @[DataMemory.scala 26:20]
  reg [31:0] ram_604; // @[DataMemory.scala 26:20]
  reg [31:0] ram_605; // @[DataMemory.scala 26:20]
  reg [31:0] ram_606; // @[DataMemory.scala 26:20]
  reg [31:0] ram_607; // @[DataMemory.scala 26:20]
  reg [31:0] ram_608; // @[DataMemory.scala 26:20]
  reg [31:0] ram_609; // @[DataMemory.scala 26:20]
  reg [31:0] ram_610; // @[DataMemory.scala 26:20]
  reg [31:0] ram_611; // @[DataMemory.scala 26:20]
  reg [31:0] ram_612; // @[DataMemory.scala 26:20]
  reg [31:0] ram_613; // @[DataMemory.scala 26:20]
  reg [31:0] ram_614; // @[DataMemory.scala 26:20]
  reg [31:0] ram_615; // @[DataMemory.scala 26:20]
  reg [31:0] ram_616; // @[DataMemory.scala 26:20]
  reg [31:0] ram_617; // @[DataMemory.scala 26:20]
  reg [31:0] ram_618; // @[DataMemory.scala 26:20]
  reg [31:0] ram_619; // @[DataMemory.scala 26:20]
  reg [31:0] ram_620; // @[DataMemory.scala 26:20]
  reg [31:0] ram_621; // @[DataMemory.scala 26:20]
  reg [31:0] ram_622; // @[DataMemory.scala 26:20]
  reg [31:0] ram_623; // @[DataMemory.scala 26:20]
  reg [31:0] ram_624; // @[DataMemory.scala 26:20]
  reg [31:0] ram_625; // @[DataMemory.scala 26:20]
  reg [31:0] ram_626; // @[DataMemory.scala 26:20]
  reg [31:0] ram_627; // @[DataMemory.scala 26:20]
  reg [31:0] ram_628; // @[DataMemory.scala 26:20]
  reg [31:0] ram_629; // @[DataMemory.scala 26:20]
  reg [31:0] ram_630; // @[DataMemory.scala 26:20]
  reg [31:0] ram_631; // @[DataMemory.scala 26:20]
  reg [31:0] ram_632; // @[DataMemory.scala 26:20]
  reg [31:0] ram_633; // @[DataMemory.scala 26:20]
  reg [31:0] ram_634; // @[DataMemory.scala 26:20]
  reg [31:0] ram_635; // @[DataMemory.scala 26:20]
  reg [31:0] ram_636; // @[DataMemory.scala 26:20]
  reg [31:0] ram_637; // @[DataMemory.scala 26:20]
  reg [31:0] ram_638; // @[DataMemory.scala 26:20]
  reg [31:0] ram_639; // @[DataMemory.scala 26:20]
  reg [31:0] ram_640; // @[DataMemory.scala 26:20]
  reg [31:0] ram_641; // @[DataMemory.scala 26:20]
  reg [31:0] ram_642; // @[DataMemory.scala 26:20]
  reg [31:0] ram_643; // @[DataMemory.scala 26:20]
  reg [31:0] ram_644; // @[DataMemory.scala 26:20]
  reg [31:0] ram_645; // @[DataMemory.scala 26:20]
  reg [31:0] ram_646; // @[DataMemory.scala 26:20]
  reg [31:0] ram_647; // @[DataMemory.scala 26:20]
  reg [31:0] ram_648; // @[DataMemory.scala 26:20]
  reg [31:0] ram_649; // @[DataMemory.scala 26:20]
  reg [31:0] ram_650; // @[DataMemory.scala 26:20]
  reg [31:0] ram_651; // @[DataMemory.scala 26:20]
  reg [31:0] ram_652; // @[DataMemory.scala 26:20]
  reg [31:0] ram_653; // @[DataMemory.scala 26:20]
  reg [31:0] ram_654; // @[DataMemory.scala 26:20]
  reg [31:0] ram_655; // @[DataMemory.scala 26:20]
  reg [31:0] ram_656; // @[DataMemory.scala 26:20]
  reg [31:0] ram_657; // @[DataMemory.scala 26:20]
  reg [31:0] ram_658; // @[DataMemory.scala 26:20]
  reg [31:0] ram_659; // @[DataMemory.scala 26:20]
  reg [31:0] ram_660; // @[DataMemory.scala 26:20]
  reg [31:0] ram_661; // @[DataMemory.scala 26:20]
  reg [31:0] ram_662; // @[DataMemory.scala 26:20]
  reg [31:0] ram_663; // @[DataMemory.scala 26:20]
  reg [31:0] ram_664; // @[DataMemory.scala 26:20]
  reg [31:0] ram_665; // @[DataMemory.scala 26:20]
  reg [31:0] ram_666; // @[DataMemory.scala 26:20]
  reg [31:0] ram_667; // @[DataMemory.scala 26:20]
  reg [31:0] ram_668; // @[DataMemory.scala 26:20]
  reg [31:0] ram_669; // @[DataMemory.scala 26:20]
  reg [31:0] ram_670; // @[DataMemory.scala 26:20]
  reg [31:0] ram_671; // @[DataMemory.scala 26:20]
  reg [31:0] ram_672; // @[DataMemory.scala 26:20]
  reg [31:0] ram_673; // @[DataMemory.scala 26:20]
  reg [31:0] ram_674; // @[DataMemory.scala 26:20]
  reg [31:0] ram_675; // @[DataMemory.scala 26:20]
  reg [31:0] ram_676; // @[DataMemory.scala 26:20]
  reg [31:0] ram_677; // @[DataMemory.scala 26:20]
  reg [31:0] ram_678; // @[DataMemory.scala 26:20]
  reg [31:0] ram_679; // @[DataMemory.scala 26:20]
  reg [31:0] ram_680; // @[DataMemory.scala 26:20]
  reg [31:0] ram_681; // @[DataMemory.scala 26:20]
  reg [31:0] ram_682; // @[DataMemory.scala 26:20]
  reg [31:0] ram_683; // @[DataMemory.scala 26:20]
  reg [31:0] ram_684; // @[DataMemory.scala 26:20]
  reg [31:0] ram_685; // @[DataMemory.scala 26:20]
  reg [31:0] ram_686; // @[DataMemory.scala 26:20]
  reg [31:0] ram_687; // @[DataMemory.scala 26:20]
  reg [31:0] ram_688; // @[DataMemory.scala 26:20]
  reg [31:0] ram_689; // @[DataMemory.scala 26:20]
  reg [31:0] ram_690; // @[DataMemory.scala 26:20]
  reg [31:0] ram_691; // @[DataMemory.scala 26:20]
  reg [31:0] ram_692; // @[DataMemory.scala 26:20]
  reg [31:0] ram_693; // @[DataMemory.scala 26:20]
  reg [31:0] ram_694; // @[DataMemory.scala 26:20]
  reg [31:0] ram_695; // @[DataMemory.scala 26:20]
  reg [31:0] ram_696; // @[DataMemory.scala 26:20]
  reg [31:0] ram_697; // @[DataMemory.scala 26:20]
  reg [31:0] ram_698; // @[DataMemory.scala 26:20]
  reg [31:0] ram_699; // @[DataMemory.scala 26:20]
  reg [31:0] ram_700; // @[DataMemory.scala 26:20]
  reg [31:0] ram_701; // @[DataMemory.scala 26:20]
  reg [31:0] ram_702; // @[DataMemory.scala 26:20]
  reg [31:0] ram_703; // @[DataMemory.scala 26:20]
  reg [31:0] ram_704; // @[DataMemory.scala 26:20]
  reg [31:0] ram_705; // @[DataMemory.scala 26:20]
  reg [31:0] ram_706; // @[DataMemory.scala 26:20]
  reg [31:0] ram_707; // @[DataMemory.scala 26:20]
  reg [31:0] ram_708; // @[DataMemory.scala 26:20]
  reg [31:0] ram_709; // @[DataMemory.scala 26:20]
  reg [31:0] ram_710; // @[DataMemory.scala 26:20]
  reg [31:0] ram_711; // @[DataMemory.scala 26:20]
  reg [31:0] ram_712; // @[DataMemory.scala 26:20]
  reg [31:0] ram_713; // @[DataMemory.scala 26:20]
  reg [31:0] ram_714; // @[DataMemory.scala 26:20]
  reg [31:0] ram_715; // @[DataMemory.scala 26:20]
  reg [31:0] ram_716; // @[DataMemory.scala 26:20]
  reg [31:0] ram_717; // @[DataMemory.scala 26:20]
  reg [31:0] ram_718; // @[DataMemory.scala 26:20]
  reg [31:0] ram_719; // @[DataMemory.scala 26:20]
  reg [31:0] ram_720; // @[DataMemory.scala 26:20]
  reg [31:0] ram_721; // @[DataMemory.scala 26:20]
  reg [31:0] ram_722; // @[DataMemory.scala 26:20]
  reg [31:0] ram_723; // @[DataMemory.scala 26:20]
  reg [31:0] ram_724; // @[DataMemory.scala 26:20]
  reg [31:0] ram_725; // @[DataMemory.scala 26:20]
  reg [31:0] ram_726; // @[DataMemory.scala 26:20]
  reg [31:0] ram_727; // @[DataMemory.scala 26:20]
  reg [31:0] ram_728; // @[DataMemory.scala 26:20]
  reg [31:0] ram_729; // @[DataMemory.scala 26:20]
  reg [31:0] ram_730; // @[DataMemory.scala 26:20]
  reg [31:0] ram_731; // @[DataMemory.scala 26:20]
  reg [31:0] ram_732; // @[DataMemory.scala 26:20]
  reg [31:0] ram_733; // @[DataMemory.scala 26:20]
  reg [31:0] ram_734; // @[DataMemory.scala 26:20]
  reg [31:0] ram_735; // @[DataMemory.scala 26:20]
  reg [31:0] ram_736; // @[DataMemory.scala 26:20]
  reg [31:0] ram_737; // @[DataMemory.scala 26:20]
  reg [31:0] ram_738; // @[DataMemory.scala 26:20]
  reg [31:0] ram_739; // @[DataMemory.scala 26:20]
  reg [31:0] ram_740; // @[DataMemory.scala 26:20]
  reg [31:0] ram_741; // @[DataMemory.scala 26:20]
  reg [31:0] ram_742; // @[DataMemory.scala 26:20]
  reg [31:0] ram_743; // @[DataMemory.scala 26:20]
  reg [31:0] ram_744; // @[DataMemory.scala 26:20]
  reg [31:0] ram_745; // @[DataMemory.scala 26:20]
  reg [31:0] ram_746; // @[DataMemory.scala 26:20]
  reg [31:0] ram_747; // @[DataMemory.scala 26:20]
  reg [31:0] ram_748; // @[DataMemory.scala 26:20]
  reg [31:0] ram_749; // @[DataMemory.scala 26:20]
  reg [31:0] ram_750; // @[DataMemory.scala 26:20]
  reg [31:0] ram_751; // @[DataMemory.scala 26:20]
  reg [31:0] ram_752; // @[DataMemory.scala 26:20]
  reg [31:0] ram_753; // @[DataMemory.scala 26:20]
  reg [31:0] ram_754; // @[DataMemory.scala 26:20]
  reg [31:0] ram_755; // @[DataMemory.scala 26:20]
  reg [31:0] ram_756; // @[DataMemory.scala 26:20]
  reg [31:0] ram_757; // @[DataMemory.scala 26:20]
  reg [31:0] ram_758; // @[DataMemory.scala 26:20]
  reg [31:0] ram_759; // @[DataMemory.scala 26:20]
  reg [31:0] ram_760; // @[DataMemory.scala 26:20]
  reg [31:0] ram_761; // @[DataMemory.scala 26:20]
  reg [31:0] ram_762; // @[DataMemory.scala 26:20]
  reg [31:0] ram_763; // @[DataMemory.scala 26:20]
  reg [31:0] ram_764; // @[DataMemory.scala 26:20]
  reg [31:0] ram_765; // @[DataMemory.scala 26:20]
  reg [31:0] ram_766; // @[DataMemory.scala 26:20]
  reg [31:0] ram_767; // @[DataMemory.scala 26:20]
  reg [31:0] ram_768; // @[DataMemory.scala 26:20]
  reg [31:0] ram_769; // @[DataMemory.scala 26:20]
  reg [31:0] ram_770; // @[DataMemory.scala 26:20]
  reg [31:0] ram_771; // @[DataMemory.scala 26:20]
  reg [31:0] ram_772; // @[DataMemory.scala 26:20]
  reg [31:0] ram_773; // @[DataMemory.scala 26:20]
  reg [31:0] ram_774; // @[DataMemory.scala 26:20]
  reg [31:0] ram_775; // @[DataMemory.scala 26:20]
  reg [31:0] ram_776; // @[DataMemory.scala 26:20]
  reg [31:0] ram_777; // @[DataMemory.scala 26:20]
  reg [31:0] ram_778; // @[DataMemory.scala 26:20]
  reg [31:0] ram_779; // @[DataMemory.scala 26:20]
  reg [31:0] ram_780; // @[DataMemory.scala 26:20]
  reg [31:0] ram_781; // @[DataMemory.scala 26:20]
  reg [31:0] ram_782; // @[DataMemory.scala 26:20]
  reg [31:0] ram_783; // @[DataMemory.scala 26:20]
  reg [31:0] ram_784; // @[DataMemory.scala 26:20]
  reg [31:0] ram_785; // @[DataMemory.scala 26:20]
  reg [31:0] ram_786; // @[DataMemory.scala 26:20]
  reg [31:0] ram_787; // @[DataMemory.scala 26:20]
  reg [31:0] ram_788; // @[DataMemory.scala 26:20]
  reg [31:0] ram_789; // @[DataMemory.scala 26:20]
  reg [31:0] ram_790; // @[DataMemory.scala 26:20]
  reg [31:0] ram_791; // @[DataMemory.scala 26:20]
  reg [31:0] ram_792; // @[DataMemory.scala 26:20]
  reg [31:0] ram_793; // @[DataMemory.scala 26:20]
  reg [31:0] ram_794; // @[DataMemory.scala 26:20]
  reg [31:0] ram_795; // @[DataMemory.scala 26:20]
  reg [31:0] ram_796; // @[DataMemory.scala 26:20]
  reg [31:0] ram_797; // @[DataMemory.scala 26:20]
  reg [31:0] ram_798; // @[DataMemory.scala 26:20]
  reg [31:0] ram_799; // @[DataMemory.scala 26:20]
  reg [31:0] ram_800; // @[DataMemory.scala 26:20]
  reg [31:0] ram_801; // @[DataMemory.scala 26:20]
  reg [31:0] ram_802; // @[DataMemory.scala 26:20]
  reg [31:0] ram_803; // @[DataMemory.scala 26:20]
  reg [31:0] ram_804; // @[DataMemory.scala 26:20]
  reg [31:0] ram_805; // @[DataMemory.scala 26:20]
  reg [31:0] ram_806; // @[DataMemory.scala 26:20]
  reg [31:0] ram_807; // @[DataMemory.scala 26:20]
  reg [31:0] ram_808; // @[DataMemory.scala 26:20]
  reg [31:0] ram_809; // @[DataMemory.scala 26:20]
  reg [31:0] ram_810; // @[DataMemory.scala 26:20]
  reg [31:0] ram_811; // @[DataMemory.scala 26:20]
  reg [31:0] ram_812; // @[DataMemory.scala 26:20]
  reg [31:0] ram_813; // @[DataMemory.scala 26:20]
  reg [31:0] ram_814; // @[DataMemory.scala 26:20]
  reg [31:0] ram_815; // @[DataMemory.scala 26:20]
  reg [31:0] ram_816; // @[DataMemory.scala 26:20]
  reg [31:0] ram_817; // @[DataMemory.scala 26:20]
  reg [31:0] ram_818; // @[DataMemory.scala 26:20]
  reg [31:0] ram_819; // @[DataMemory.scala 26:20]
  reg [31:0] ram_820; // @[DataMemory.scala 26:20]
  reg [31:0] ram_821; // @[DataMemory.scala 26:20]
  reg [31:0] ram_822; // @[DataMemory.scala 26:20]
  reg [31:0] ram_823; // @[DataMemory.scala 26:20]
  reg [31:0] ram_824; // @[DataMemory.scala 26:20]
  reg [31:0] ram_825; // @[DataMemory.scala 26:20]
  reg [31:0] ram_826; // @[DataMemory.scala 26:20]
  reg [31:0] ram_827; // @[DataMemory.scala 26:20]
  reg [31:0] ram_828; // @[DataMemory.scala 26:20]
  reg [31:0] ram_829; // @[DataMemory.scala 26:20]
  reg [31:0] ram_830; // @[DataMemory.scala 26:20]
  reg [31:0] ram_831; // @[DataMemory.scala 26:20]
  reg [31:0] ram_832; // @[DataMemory.scala 26:20]
  reg [31:0] ram_833; // @[DataMemory.scala 26:20]
  reg [31:0] ram_834; // @[DataMemory.scala 26:20]
  reg [31:0] ram_835; // @[DataMemory.scala 26:20]
  reg [31:0] ram_836; // @[DataMemory.scala 26:20]
  reg [31:0] ram_837; // @[DataMemory.scala 26:20]
  reg [31:0] ram_838; // @[DataMemory.scala 26:20]
  reg [31:0] ram_839; // @[DataMemory.scala 26:20]
  reg [31:0] ram_840; // @[DataMemory.scala 26:20]
  reg [31:0] ram_841; // @[DataMemory.scala 26:20]
  reg [31:0] ram_842; // @[DataMemory.scala 26:20]
  reg [31:0] ram_843; // @[DataMemory.scala 26:20]
  reg [31:0] ram_844; // @[DataMemory.scala 26:20]
  reg [31:0] ram_845; // @[DataMemory.scala 26:20]
  reg [31:0] ram_846; // @[DataMemory.scala 26:20]
  reg [31:0] ram_847; // @[DataMemory.scala 26:20]
  reg [31:0] ram_848; // @[DataMemory.scala 26:20]
  reg [31:0] ram_849; // @[DataMemory.scala 26:20]
  reg [31:0] ram_850; // @[DataMemory.scala 26:20]
  reg [31:0] ram_851; // @[DataMemory.scala 26:20]
  reg [31:0] ram_852; // @[DataMemory.scala 26:20]
  reg [31:0] ram_853; // @[DataMemory.scala 26:20]
  reg [31:0] ram_854; // @[DataMemory.scala 26:20]
  reg [31:0] ram_855; // @[DataMemory.scala 26:20]
  reg [31:0] ram_856; // @[DataMemory.scala 26:20]
  reg [31:0] ram_857; // @[DataMemory.scala 26:20]
  reg [31:0] ram_858; // @[DataMemory.scala 26:20]
  reg [31:0] ram_859; // @[DataMemory.scala 26:20]
  reg [31:0] ram_860; // @[DataMemory.scala 26:20]
  reg [31:0] ram_861; // @[DataMemory.scala 26:20]
  reg [31:0] ram_862; // @[DataMemory.scala 26:20]
  reg [31:0] ram_863; // @[DataMemory.scala 26:20]
  reg [31:0] ram_864; // @[DataMemory.scala 26:20]
  reg [31:0] ram_865; // @[DataMemory.scala 26:20]
  reg [31:0] ram_866; // @[DataMemory.scala 26:20]
  reg [31:0] ram_867; // @[DataMemory.scala 26:20]
  reg [31:0] ram_868; // @[DataMemory.scala 26:20]
  reg [31:0] ram_869; // @[DataMemory.scala 26:20]
  reg [31:0] ram_870; // @[DataMemory.scala 26:20]
  reg [31:0] ram_871; // @[DataMemory.scala 26:20]
  reg [31:0] ram_872; // @[DataMemory.scala 26:20]
  reg [31:0] ram_873; // @[DataMemory.scala 26:20]
  reg [31:0] ram_874; // @[DataMemory.scala 26:20]
  reg [31:0] ram_875; // @[DataMemory.scala 26:20]
  reg [31:0] ram_876; // @[DataMemory.scala 26:20]
  reg [31:0] ram_877; // @[DataMemory.scala 26:20]
  reg [31:0] ram_878; // @[DataMemory.scala 26:20]
  reg [31:0] ram_879; // @[DataMemory.scala 26:20]
  reg [31:0] ram_880; // @[DataMemory.scala 26:20]
  reg [31:0] ram_881; // @[DataMemory.scala 26:20]
  reg [31:0] ram_882; // @[DataMemory.scala 26:20]
  reg [31:0] ram_883; // @[DataMemory.scala 26:20]
  reg [31:0] ram_884; // @[DataMemory.scala 26:20]
  reg [31:0] ram_885; // @[DataMemory.scala 26:20]
  reg [31:0] ram_886; // @[DataMemory.scala 26:20]
  reg [31:0] ram_887; // @[DataMemory.scala 26:20]
  reg [31:0] ram_888; // @[DataMemory.scala 26:20]
  reg [31:0] ram_889; // @[DataMemory.scala 26:20]
  reg [31:0] ram_890; // @[DataMemory.scala 26:20]
  reg [31:0] ram_891; // @[DataMemory.scala 26:20]
  reg [31:0] ram_892; // @[DataMemory.scala 26:20]
  reg [31:0] ram_893; // @[DataMemory.scala 26:20]
  reg [31:0] ram_894; // @[DataMemory.scala 26:20]
  reg [31:0] ram_895; // @[DataMemory.scala 26:20]
  reg [31:0] ram_896; // @[DataMemory.scala 26:20]
  reg [31:0] ram_897; // @[DataMemory.scala 26:20]
  reg [31:0] ram_898; // @[DataMemory.scala 26:20]
  reg [31:0] ram_899; // @[DataMemory.scala 26:20]
  reg [31:0] ram_900; // @[DataMemory.scala 26:20]
  reg [31:0] ram_901; // @[DataMemory.scala 26:20]
  reg [31:0] ram_902; // @[DataMemory.scala 26:20]
  reg [31:0] ram_903; // @[DataMemory.scala 26:20]
  reg [31:0] ram_904; // @[DataMemory.scala 26:20]
  reg [31:0] ram_905; // @[DataMemory.scala 26:20]
  reg [31:0] ram_906; // @[DataMemory.scala 26:20]
  reg [31:0] ram_907; // @[DataMemory.scala 26:20]
  reg [31:0] ram_908; // @[DataMemory.scala 26:20]
  reg [31:0] ram_909; // @[DataMemory.scala 26:20]
  reg [31:0] ram_910; // @[DataMemory.scala 26:20]
  reg [31:0] ram_911; // @[DataMemory.scala 26:20]
  reg [31:0] ram_912; // @[DataMemory.scala 26:20]
  reg [31:0] ram_913; // @[DataMemory.scala 26:20]
  reg [31:0] ram_914; // @[DataMemory.scala 26:20]
  reg [31:0] ram_915; // @[DataMemory.scala 26:20]
  reg [31:0] ram_916; // @[DataMemory.scala 26:20]
  reg [31:0] ram_917; // @[DataMemory.scala 26:20]
  reg [31:0] ram_918; // @[DataMemory.scala 26:20]
  reg [31:0] ram_919; // @[DataMemory.scala 26:20]
  reg [31:0] ram_920; // @[DataMemory.scala 26:20]
  reg [31:0] ram_921; // @[DataMemory.scala 26:20]
  reg [31:0] ram_922; // @[DataMemory.scala 26:20]
  reg [31:0] ram_923; // @[DataMemory.scala 26:20]
  reg [31:0] ram_924; // @[DataMemory.scala 26:20]
  reg [31:0] ram_925; // @[DataMemory.scala 26:20]
  reg [31:0] ram_926; // @[DataMemory.scala 26:20]
  reg [31:0] ram_927; // @[DataMemory.scala 26:20]
  reg [31:0] ram_928; // @[DataMemory.scala 26:20]
  reg [31:0] ram_929; // @[DataMemory.scala 26:20]
  reg [31:0] ram_930; // @[DataMemory.scala 26:20]
  reg [31:0] ram_931; // @[DataMemory.scala 26:20]
  reg [31:0] ram_932; // @[DataMemory.scala 26:20]
  reg [31:0] ram_933; // @[DataMemory.scala 26:20]
  reg [31:0] ram_934; // @[DataMemory.scala 26:20]
  reg [31:0] ram_935; // @[DataMemory.scala 26:20]
  reg [31:0] ram_936; // @[DataMemory.scala 26:20]
  reg [31:0] ram_937; // @[DataMemory.scala 26:20]
  reg [31:0] ram_938; // @[DataMemory.scala 26:20]
  reg [31:0] ram_939; // @[DataMemory.scala 26:20]
  reg [31:0] ram_940; // @[DataMemory.scala 26:20]
  reg [31:0] ram_941; // @[DataMemory.scala 26:20]
  reg [31:0] ram_942; // @[DataMemory.scala 26:20]
  reg [31:0] ram_943; // @[DataMemory.scala 26:20]
  reg [31:0] ram_944; // @[DataMemory.scala 26:20]
  reg [31:0] ram_945; // @[DataMemory.scala 26:20]
  reg [31:0] ram_946; // @[DataMemory.scala 26:20]
  reg [31:0] ram_947; // @[DataMemory.scala 26:20]
  reg [31:0] ram_948; // @[DataMemory.scala 26:20]
  reg [31:0] ram_949; // @[DataMemory.scala 26:20]
  reg [31:0] ram_950; // @[DataMemory.scala 26:20]
  reg [31:0] ram_951; // @[DataMemory.scala 26:20]
  reg [31:0] ram_952; // @[DataMemory.scala 26:20]
  reg [31:0] ram_953; // @[DataMemory.scala 26:20]
  reg [31:0] ram_954; // @[DataMemory.scala 26:20]
  reg [31:0] ram_955; // @[DataMemory.scala 26:20]
  reg [31:0] ram_956; // @[DataMemory.scala 26:20]
  reg [31:0] ram_957; // @[DataMemory.scala 26:20]
  reg [31:0] ram_958; // @[DataMemory.scala 26:20]
  reg [31:0] ram_959; // @[DataMemory.scala 26:20]
  reg [31:0] ram_960; // @[DataMemory.scala 26:20]
  reg [31:0] ram_961; // @[DataMemory.scala 26:20]
  reg [31:0] ram_962; // @[DataMemory.scala 26:20]
  reg [31:0] ram_963; // @[DataMemory.scala 26:20]
  reg [31:0] ram_964; // @[DataMemory.scala 26:20]
  reg [31:0] ram_965; // @[DataMemory.scala 26:20]
  reg [31:0] ram_966; // @[DataMemory.scala 26:20]
  reg [31:0] ram_967; // @[DataMemory.scala 26:20]
  reg [31:0] ram_968; // @[DataMemory.scala 26:20]
  reg [31:0] ram_969; // @[DataMemory.scala 26:20]
  reg [31:0] ram_970; // @[DataMemory.scala 26:20]
  reg [31:0] ram_971; // @[DataMemory.scala 26:20]
  reg [31:0] ram_972; // @[DataMemory.scala 26:20]
  reg [31:0] ram_973; // @[DataMemory.scala 26:20]
  reg [31:0] ram_974; // @[DataMemory.scala 26:20]
  reg [31:0] ram_975; // @[DataMemory.scala 26:20]
  reg [31:0] ram_976; // @[DataMemory.scala 26:20]
  reg [31:0] ram_977; // @[DataMemory.scala 26:20]
  reg [31:0] ram_978; // @[DataMemory.scala 26:20]
  reg [31:0] ram_979; // @[DataMemory.scala 26:20]
  reg [31:0] ram_980; // @[DataMemory.scala 26:20]
  reg [31:0] ram_981; // @[DataMemory.scala 26:20]
  reg [31:0] ram_982; // @[DataMemory.scala 26:20]
  reg [31:0] ram_983; // @[DataMemory.scala 26:20]
  reg [31:0] ram_984; // @[DataMemory.scala 26:20]
  reg [31:0] ram_985; // @[DataMemory.scala 26:20]
  reg [31:0] ram_986; // @[DataMemory.scala 26:20]
  reg [31:0] ram_987; // @[DataMemory.scala 26:20]
  reg [31:0] ram_988; // @[DataMemory.scala 26:20]
  reg [31:0] ram_989; // @[DataMemory.scala 26:20]
  reg [31:0] ram_990; // @[DataMemory.scala 26:20]
  reg [31:0] ram_991; // @[DataMemory.scala 26:20]
  reg [31:0] ram_992; // @[DataMemory.scala 26:20]
  reg [31:0] ram_993; // @[DataMemory.scala 26:20]
  reg [31:0] ram_994; // @[DataMemory.scala 26:20]
  reg [31:0] ram_995; // @[DataMemory.scala 26:20]
  reg [31:0] ram_996; // @[DataMemory.scala 26:20]
  reg [31:0] ram_997; // @[DataMemory.scala 26:20]
  reg [31:0] ram_998; // @[DataMemory.scala 26:20]
  reg [31:0] ram_999; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1000; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1001; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1002; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1003; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1004; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1005; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1006; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1007; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1008; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1009; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1010; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1011; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1012; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1013; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1014; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1015; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1016; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1017; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1018; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1019; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1020; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1021; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1022; // @[DataMemory.scala 26:20]
  reg [31:0] ram_1023; // @[DataMemory.scala 26:20]
  wire [31:0] _GEN_1 = 8'h1 == io_addr[9:2] ? ram_1 : ram_0; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_2 = 8'h2 == io_addr[9:2] ? ram_2 : _GEN_1; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_3 = 8'h3 == io_addr[9:2] ? ram_3 : _GEN_2; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_4 = 8'h4 == io_addr[9:2] ? ram_4 : _GEN_3; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_5 = 8'h5 == io_addr[9:2] ? ram_5 : _GEN_4; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_6 = 8'h6 == io_addr[9:2] ? ram_6 : _GEN_5; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_7 = 8'h7 == io_addr[9:2] ? ram_7 : _GEN_6; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_8 = 8'h8 == io_addr[9:2] ? ram_8 : _GEN_7; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_9 = 8'h9 == io_addr[9:2] ? ram_9 : _GEN_8; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_10 = 8'ha == io_addr[9:2] ? ram_10 : _GEN_9; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_11 = 8'hb == io_addr[9:2] ? ram_11 : _GEN_10; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_12 = 8'hc == io_addr[9:2] ? ram_12 : _GEN_11; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_13 = 8'hd == io_addr[9:2] ? ram_13 : _GEN_12; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_14 = 8'he == io_addr[9:2] ? ram_14 : _GEN_13; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_15 = 8'hf == io_addr[9:2] ? ram_15 : _GEN_14; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_16 = 8'h10 == io_addr[9:2] ? ram_16 : _GEN_15; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_17 = 8'h11 == io_addr[9:2] ? ram_17 : _GEN_16; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_18 = 8'h12 == io_addr[9:2] ? ram_18 : _GEN_17; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_19 = 8'h13 == io_addr[9:2] ? ram_19 : _GEN_18; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_20 = 8'h14 == io_addr[9:2] ? ram_20 : _GEN_19; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_21 = 8'h15 == io_addr[9:2] ? ram_21 : _GEN_20; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_22 = 8'h16 == io_addr[9:2] ? ram_22 : _GEN_21; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_23 = 8'h17 == io_addr[9:2] ? ram_23 : _GEN_22; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_24 = 8'h18 == io_addr[9:2] ? ram_24 : _GEN_23; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_25 = 8'h19 == io_addr[9:2] ? ram_25 : _GEN_24; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_26 = 8'h1a == io_addr[9:2] ? ram_26 : _GEN_25; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_27 = 8'h1b == io_addr[9:2] ? ram_27 : _GEN_26; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_28 = 8'h1c == io_addr[9:2] ? ram_28 : _GEN_27; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_29 = 8'h1d == io_addr[9:2] ? ram_29 : _GEN_28; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_30 = 8'h1e == io_addr[9:2] ? ram_30 : _GEN_29; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_31 = 8'h1f == io_addr[9:2] ? ram_31 : _GEN_30; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_32 = 8'h20 == io_addr[9:2] ? ram_32 : _GEN_31; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_33 = 8'h21 == io_addr[9:2] ? ram_33 : _GEN_32; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_34 = 8'h22 == io_addr[9:2] ? ram_34 : _GEN_33; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_35 = 8'h23 == io_addr[9:2] ? ram_35 : _GEN_34; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_36 = 8'h24 == io_addr[9:2] ? ram_36 : _GEN_35; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_37 = 8'h25 == io_addr[9:2] ? ram_37 : _GEN_36; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_38 = 8'h26 == io_addr[9:2] ? ram_38 : _GEN_37; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_39 = 8'h27 == io_addr[9:2] ? ram_39 : _GEN_38; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_40 = 8'h28 == io_addr[9:2] ? ram_40 : _GEN_39; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_41 = 8'h29 == io_addr[9:2] ? ram_41 : _GEN_40; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_42 = 8'h2a == io_addr[9:2] ? ram_42 : _GEN_41; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_43 = 8'h2b == io_addr[9:2] ? ram_43 : _GEN_42; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_44 = 8'h2c == io_addr[9:2] ? ram_44 : _GEN_43; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_45 = 8'h2d == io_addr[9:2] ? ram_45 : _GEN_44; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_46 = 8'h2e == io_addr[9:2] ? ram_46 : _GEN_45; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_47 = 8'h2f == io_addr[9:2] ? ram_47 : _GEN_46; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_48 = 8'h30 == io_addr[9:2] ? ram_48 : _GEN_47; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_49 = 8'h31 == io_addr[9:2] ? ram_49 : _GEN_48; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_50 = 8'h32 == io_addr[9:2] ? ram_50 : _GEN_49; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_51 = 8'h33 == io_addr[9:2] ? ram_51 : _GEN_50; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_52 = 8'h34 == io_addr[9:2] ? ram_52 : _GEN_51; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_53 = 8'h35 == io_addr[9:2] ? ram_53 : _GEN_52; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_54 = 8'h36 == io_addr[9:2] ? ram_54 : _GEN_53; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_55 = 8'h37 == io_addr[9:2] ? ram_55 : _GEN_54; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_56 = 8'h38 == io_addr[9:2] ? ram_56 : _GEN_55; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_57 = 8'h39 == io_addr[9:2] ? ram_57 : _GEN_56; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_58 = 8'h3a == io_addr[9:2] ? ram_58 : _GEN_57; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_59 = 8'h3b == io_addr[9:2] ? ram_59 : _GEN_58; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_60 = 8'h3c == io_addr[9:2] ? ram_60 : _GEN_59; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_61 = 8'h3d == io_addr[9:2] ? ram_61 : _GEN_60; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_62 = 8'h3e == io_addr[9:2] ? ram_62 : _GEN_61; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_63 = 8'h3f == io_addr[9:2] ? ram_63 : _GEN_62; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_64 = 8'h40 == io_addr[9:2] ? ram_64 : _GEN_63; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_65 = 8'h41 == io_addr[9:2] ? ram_65 : _GEN_64; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_66 = 8'h42 == io_addr[9:2] ? ram_66 : _GEN_65; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_67 = 8'h43 == io_addr[9:2] ? ram_67 : _GEN_66; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_68 = 8'h44 == io_addr[9:2] ? ram_68 : _GEN_67; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_69 = 8'h45 == io_addr[9:2] ? ram_69 : _GEN_68; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_70 = 8'h46 == io_addr[9:2] ? ram_70 : _GEN_69; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_71 = 8'h47 == io_addr[9:2] ? ram_71 : _GEN_70; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_72 = 8'h48 == io_addr[9:2] ? ram_72 : _GEN_71; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_73 = 8'h49 == io_addr[9:2] ? ram_73 : _GEN_72; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_74 = 8'h4a == io_addr[9:2] ? ram_74 : _GEN_73; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_75 = 8'h4b == io_addr[9:2] ? ram_75 : _GEN_74; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_76 = 8'h4c == io_addr[9:2] ? ram_76 : _GEN_75; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_77 = 8'h4d == io_addr[9:2] ? ram_77 : _GEN_76; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_78 = 8'h4e == io_addr[9:2] ? ram_78 : _GEN_77; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_79 = 8'h4f == io_addr[9:2] ? ram_79 : _GEN_78; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_80 = 8'h50 == io_addr[9:2] ? ram_80 : _GEN_79; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_81 = 8'h51 == io_addr[9:2] ? ram_81 : _GEN_80; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_82 = 8'h52 == io_addr[9:2] ? ram_82 : _GEN_81; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_83 = 8'h53 == io_addr[9:2] ? ram_83 : _GEN_82; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_84 = 8'h54 == io_addr[9:2] ? ram_84 : _GEN_83; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_85 = 8'h55 == io_addr[9:2] ? ram_85 : _GEN_84; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_86 = 8'h56 == io_addr[9:2] ? ram_86 : _GEN_85; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_87 = 8'h57 == io_addr[9:2] ? ram_87 : _GEN_86; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_88 = 8'h58 == io_addr[9:2] ? ram_88 : _GEN_87; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_89 = 8'h59 == io_addr[9:2] ? ram_89 : _GEN_88; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_90 = 8'h5a == io_addr[9:2] ? ram_90 : _GEN_89; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_91 = 8'h5b == io_addr[9:2] ? ram_91 : _GEN_90; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_92 = 8'h5c == io_addr[9:2] ? ram_92 : _GEN_91; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_93 = 8'h5d == io_addr[9:2] ? ram_93 : _GEN_92; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_94 = 8'h5e == io_addr[9:2] ? ram_94 : _GEN_93; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_95 = 8'h5f == io_addr[9:2] ? ram_95 : _GEN_94; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_96 = 8'h60 == io_addr[9:2] ? ram_96 : _GEN_95; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_97 = 8'h61 == io_addr[9:2] ? ram_97 : _GEN_96; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_98 = 8'h62 == io_addr[9:2] ? ram_98 : _GEN_97; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_99 = 8'h63 == io_addr[9:2] ? ram_99 : _GEN_98; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_100 = 8'h64 == io_addr[9:2] ? ram_100 : _GEN_99; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_101 = 8'h65 == io_addr[9:2] ? ram_101 : _GEN_100; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_102 = 8'h66 == io_addr[9:2] ? ram_102 : _GEN_101; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_103 = 8'h67 == io_addr[9:2] ? ram_103 : _GEN_102; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_104 = 8'h68 == io_addr[9:2] ? ram_104 : _GEN_103; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_105 = 8'h69 == io_addr[9:2] ? ram_105 : _GEN_104; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_106 = 8'h6a == io_addr[9:2] ? ram_106 : _GEN_105; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_107 = 8'h6b == io_addr[9:2] ? ram_107 : _GEN_106; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_108 = 8'h6c == io_addr[9:2] ? ram_108 : _GEN_107; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_109 = 8'h6d == io_addr[9:2] ? ram_109 : _GEN_108; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_110 = 8'h6e == io_addr[9:2] ? ram_110 : _GEN_109; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_111 = 8'h6f == io_addr[9:2] ? ram_111 : _GEN_110; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_112 = 8'h70 == io_addr[9:2] ? ram_112 : _GEN_111; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_113 = 8'h71 == io_addr[9:2] ? ram_113 : _GEN_112; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_114 = 8'h72 == io_addr[9:2] ? ram_114 : _GEN_113; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_115 = 8'h73 == io_addr[9:2] ? ram_115 : _GEN_114; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_116 = 8'h74 == io_addr[9:2] ? ram_116 : _GEN_115; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_117 = 8'h75 == io_addr[9:2] ? ram_117 : _GEN_116; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_118 = 8'h76 == io_addr[9:2] ? ram_118 : _GEN_117; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_119 = 8'h77 == io_addr[9:2] ? ram_119 : _GEN_118; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_120 = 8'h78 == io_addr[9:2] ? ram_120 : _GEN_119; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_121 = 8'h79 == io_addr[9:2] ? ram_121 : _GEN_120; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_122 = 8'h7a == io_addr[9:2] ? ram_122 : _GEN_121; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_123 = 8'h7b == io_addr[9:2] ? ram_123 : _GEN_122; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_124 = 8'h7c == io_addr[9:2] ? ram_124 : _GEN_123; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_125 = 8'h7d == io_addr[9:2] ? ram_125 : _GEN_124; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_126 = 8'h7e == io_addr[9:2] ? ram_126 : _GEN_125; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_127 = 8'h7f == io_addr[9:2] ? ram_127 : _GEN_126; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_128 = 8'h80 == io_addr[9:2] ? ram_128 : _GEN_127; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_129 = 8'h81 == io_addr[9:2] ? ram_129 : _GEN_128; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_130 = 8'h82 == io_addr[9:2] ? ram_130 : _GEN_129; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_131 = 8'h83 == io_addr[9:2] ? ram_131 : _GEN_130; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_132 = 8'h84 == io_addr[9:2] ? ram_132 : _GEN_131; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_133 = 8'h85 == io_addr[9:2] ? ram_133 : _GEN_132; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_134 = 8'h86 == io_addr[9:2] ? ram_134 : _GEN_133; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_135 = 8'h87 == io_addr[9:2] ? ram_135 : _GEN_134; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_136 = 8'h88 == io_addr[9:2] ? ram_136 : _GEN_135; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_137 = 8'h89 == io_addr[9:2] ? ram_137 : _GEN_136; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_138 = 8'h8a == io_addr[9:2] ? ram_138 : _GEN_137; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_139 = 8'h8b == io_addr[9:2] ? ram_139 : _GEN_138; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_140 = 8'h8c == io_addr[9:2] ? ram_140 : _GEN_139; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_141 = 8'h8d == io_addr[9:2] ? ram_141 : _GEN_140; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_142 = 8'h8e == io_addr[9:2] ? ram_142 : _GEN_141; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_143 = 8'h8f == io_addr[9:2] ? ram_143 : _GEN_142; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_144 = 8'h90 == io_addr[9:2] ? ram_144 : _GEN_143; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_145 = 8'h91 == io_addr[9:2] ? ram_145 : _GEN_144; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_146 = 8'h92 == io_addr[9:2] ? ram_146 : _GEN_145; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_147 = 8'h93 == io_addr[9:2] ? ram_147 : _GEN_146; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_148 = 8'h94 == io_addr[9:2] ? ram_148 : _GEN_147; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_149 = 8'h95 == io_addr[9:2] ? ram_149 : _GEN_148; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_150 = 8'h96 == io_addr[9:2] ? ram_150 : _GEN_149; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_151 = 8'h97 == io_addr[9:2] ? ram_151 : _GEN_150; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_152 = 8'h98 == io_addr[9:2] ? ram_152 : _GEN_151; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_153 = 8'h99 == io_addr[9:2] ? ram_153 : _GEN_152; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_154 = 8'h9a == io_addr[9:2] ? ram_154 : _GEN_153; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_155 = 8'h9b == io_addr[9:2] ? ram_155 : _GEN_154; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_156 = 8'h9c == io_addr[9:2] ? ram_156 : _GEN_155; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_157 = 8'h9d == io_addr[9:2] ? ram_157 : _GEN_156; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_158 = 8'h9e == io_addr[9:2] ? ram_158 : _GEN_157; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_159 = 8'h9f == io_addr[9:2] ? ram_159 : _GEN_158; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_160 = 8'ha0 == io_addr[9:2] ? ram_160 : _GEN_159; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_161 = 8'ha1 == io_addr[9:2] ? ram_161 : _GEN_160; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_162 = 8'ha2 == io_addr[9:2] ? ram_162 : _GEN_161; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_163 = 8'ha3 == io_addr[9:2] ? ram_163 : _GEN_162; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_164 = 8'ha4 == io_addr[9:2] ? ram_164 : _GEN_163; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_165 = 8'ha5 == io_addr[9:2] ? ram_165 : _GEN_164; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_166 = 8'ha6 == io_addr[9:2] ? ram_166 : _GEN_165; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_167 = 8'ha7 == io_addr[9:2] ? ram_167 : _GEN_166; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_168 = 8'ha8 == io_addr[9:2] ? ram_168 : _GEN_167; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_169 = 8'ha9 == io_addr[9:2] ? ram_169 : _GEN_168; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_170 = 8'haa == io_addr[9:2] ? ram_170 : _GEN_169; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_171 = 8'hab == io_addr[9:2] ? ram_171 : _GEN_170; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_172 = 8'hac == io_addr[9:2] ? ram_172 : _GEN_171; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_173 = 8'had == io_addr[9:2] ? ram_173 : _GEN_172; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_174 = 8'hae == io_addr[9:2] ? ram_174 : _GEN_173; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_175 = 8'haf == io_addr[9:2] ? ram_175 : _GEN_174; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_176 = 8'hb0 == io_addr[9:2] ? ram_176 : _GEN_175; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_177 = 8'hb1 == io_addr[9:2] ? ram_177 : _GEN_176; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_178 = 8'hb2 == io_addr[9:2] ? ram_178 : _GEN_177; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_179 = 8'hb3 == io_addr[9:2] ? ram_179 : _GEN_178; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_180 = 8'hb4 == io_addr[9:2] ? ram_180 : _GEN_179; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_181 = 8'hb5 == io_addr[9:2] ? ram_181 : _GEN_180; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_182 = 8'hb6 == io_addr[9:2] ? ram_182 : _GEN_181; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_183 = 8'hb7 == io_addr[9:2] ? ram_183 : _GEN_182; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_184 = 8'hb8 == io_addr[9:2] ? ram_184 : _GEN_183; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_185 = 8'hb9 == io_addr[9:2] ? ram_185 : _GEN_184; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_186 = 8'hba == io_addr[9:2] ? ram_186 : _GEN_185; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_187 = 8'hbb == io_addr[9:2] ? ram_187 : _GEN_186; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_188 = 8'hbc == io_addr[9:2] ? ram_188 : _GEN_187; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_189 = 8'hbd == io_addr[9:2] ? ram_189 : _GEN_188; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_190 = 8'hbe == io_addr[9:2] ? ram_190 : _GEN_189; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_191 = 8'hbf == io_addr[9:2] ? ram_191 : _GEN_190; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_192 = 8'hc0 == io_addr[9:2] ? ram_192 : _GEN_191; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_193 = 8'hc1 == io_addr[9:2] ? ram_193 : _GEN_192; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_194 = 8'hc2 == io_addr[9:2] ? ram_194 : _GEN_193; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_195 = 8'hc3 == io_addr[9:2] ? ram_195 : _GEN_194; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_196 = 8'hc4 == io_addr[9:2] ? ram_196 : _GEN_195; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_197 = 8'hc5 == io_addr[9:2] ? ram_197 : _GEN_196; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_198 = 8'hc6 == io_addr[9:2] ? ram_198 : _GEN_197; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_199 = 8'hc7 == io_addr[9:2] ? ram_199 : _GEN_198; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_200 = 8'hc8 == io_addr[9:2] ? ram_200 : _GEN_199; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_201 = 8'hc9 == io_addr[9:2] ? ram_201 : _GEN_200; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_202 = 8'hca == io_addr[9:2] ? ram_202 : _GEN_201; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_203 = 8'hcb == io_addr[9:2] ? ram_203 : _GEN_202; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_204 = 8'hcc == io_addr[9:2] ? ram_204 : _GEN_203; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_205 = 8'hcd == io_addr[9:2] ? ram_205 : _GEN_204; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_206 = 8'hce == io_addr[9:2] ? ram_206 : _GEN_205; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_207 = 8'hcf == io_addr[9:2] ? ram_207 : _GEN_206; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_208 = 8'hd0 == io_addr[9:2] ? ram_208 : _GEN_207; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_209 = 8'hd1 == io_addr[9:2] ? ram_209 : _GEN_208; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_210 = 8'hd2 == io_addr[9:2] ? ram_210 : _GEN_209; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_211 = 8'hd3 == io_addr[9:2] ? ram_211 : _GEN_210; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_212 = 8'hd4 == io_addr[9:2] ? ram_212 : _GEN_211; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_213 = 8'hd5 == io_addr[9:2] ? ram_213 : _GEN_212; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_214 = 8'hd6 == io_addr[9:2] ? ram_214 : _GEN_213; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_215 = 8'hd7 == io_addr[9:2] ? ram_215 : _GEN_214; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_216 = 8'hd8 == io_addr[9:2] ? ram_216 : _GEN_215; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_217 = 8'hd9 == io_addr[9:2] ? ram_217 : _GEN_216; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_218 = 8'hda == io_addr[9:2] ? ram_218 : _GEN_217; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_219 = 8'hdb == io_addr[9:2] ? ram_219 : _GEN_218; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_220 = 8'hdc == io_addr[9:2] ? ram_220 : _GEN_219; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_221 = 8'hdd == io_addr[9:2] ? ram_221 : _GEN_220; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_222 = 8'hde == io_addr[9:2] ? ram_222 : _GEN_221; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_223 = 8'hdf == io_addr[9:2] ? ram_223 : _GEN_222; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_224 = 8'he0 == io_addr[9:2] ? ram_224 : _GEN_223; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_225 = 8'he1 == io_addr[9:2] ? ram_225 : _GEN_224; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_226 = 8'he2 == io_addr[9:2] ? ram_226 : _GEN_225; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_227 = 8'he3 == io_addr[9:2] ? ram_227 : _GEN_226; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_228 = 8'he4 == io_addr[9:2] ? ram_228 : _GEN_227; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_229 = 8'he5 == io_addr[9:2] ? ram_229 : _GEN_228; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_230 = 8'he6 == io_addr[9:2] ? ram_230 : _GEN_229; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_231 = 8'he7 == io_addr[9:2] ? ram_231 : _GEN_230; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_232 = 8'he8 == io_addr[9:2] ? ram_232 : _GEN_231; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_233 = 8'he9 == io_addr[9:2] ? ram_233 : _GEN_232; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_234 = 8'hea == io_addr[9:2] ? ram_234 : _GEN_233; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_235 = 8'heb == io_addr[9:2] ? ram_235 : _GEN_234; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_236 = 8'hec == io_addr[9:2] ? ram_236 : _GEN_235; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_237 = 8'hed == io_addr[9:2] ? ram_237 : _GEN_236; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_238 = 8'hee == io_addr[9:2] ? ram_238 : _GEN_237; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_239 = 8'hef == io_addr[9:2] ? ram_239 : _GEN_238; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_240 = 8'hf0 == io_addr[9:2] ? ram_240 : _GEN_239; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_241 = 8'hf1 == io_addr[9:2] ? ram_241 : _GEN_240; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_242 = 8'hf2 == io_addr[9:2] ? ram_242 : _GEN_241; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_243 = 8'hf3 == io_addr[9:2] ? ram_243 : _GEN_242; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_244 = 8'hf4 == io_addr[9:2] ? ram_244 : _GEN_243; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_245 = 8'hf5 == io_addr[9:2] ? ram_245 : _GEN_244; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_246 = 8'hf6 == io_addr[9:2] ? ram_246 : _GEN_245; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_247 = 8'hf7 == io_addr[9:2] ? ram_247 : _GEN_246; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_248 = 8'hf8 == io_addr[9:2] ? ram_248 : _GEN_247; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_249 = 8'hf9 == io_addr[9:2] ? ram_249 : _GEN_248; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_250 = 8'hfa == io_addr[9:2] ? ram_250 : _GEN_249; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_251 = 8'hfb == io_addr[9:2] ? ram_251 : _GEN_250; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_252 = 8'hfc == io_addr[9:2] ? ram_252 : _GEN_251; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_253 = 8'hfd == io_addr[9:2] ? ram_253 : _GEN_252; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_254 = 8'hfe == io_addr[9:2] ? ram_254 : _GEN_253; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_255 = 8'hff == io_addr[9:2] ? ram_255 : _GEN_254; // @[DataMemory.scala 42:{28,28}]
  wire [8:0] _GEN_7170 = {{1'd0}, io_addr[9:2]}; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_256 = 9'h100 == _GEN_7170 ? ram_256 : _GEN_255; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_257 = 9'h101 == _GEN_7170 ? ram_257 : _GEN_256; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_258 = 9'h102 == _GEN_7170 ? ram_258 : _GEN_257; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_259 = 9'h103 == _GEN_7170 ? ram_259 : _GEN_258; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_260 = 9'h104 == _GEN_7170 ? ram_260 : _GEN_259; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_261 = 9'h105 == _GEN_7170 ? ram_261 : _GEN_260; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_262 = 9'h106 == _GEN_7170 ? ram_262 : _GEN_261; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_263 = 9'h107 == _GEN_7170 ? ram_263 : _GEN_262; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_264 = 9'h108 == _GEN_7170 ? ram_264 : _GEN_263; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_265 = 9'h109 == _GEN_7170 ? ram_265 : _GEN_264; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_266 = 9'h10a == _GEN_7170 ? ram_266 : _GEN_265; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_267 = 9'h10b == _GEN_7170 ? ram_267 : _GEN_266; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_268 = 9'h10c == _GEN_7170 ? ram_268 : _GEN_267; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_269 = 9'h10d == _GEN_7170 ? ram_269 : _GEN_268; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_270 = 9'h10e == _GEN_7170 ? ram_270 : _GEN_269; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_271 = 9'h10f == _GEN_7170 ? ram_271 : _GEN_270; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_272 = 9'h110 == _GEN_7170 ? ram_272 : _GEN_271; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_273 = 9'h111 == _GEN_7170 ? ram_273 : _GEN_272; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_274 = 9'h112 == _GEN_7170 ? ram_274 : _GEN_273; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_275 = 9'h113 == _GEN_7170 ? ram_275 : _GEN_274; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_276 = 9'h114 == _GEN_7170 ? ram_276 : _GEN_275; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_277 = 9'h115 == _GEN_7170 ? ram_277 : _GEN_276; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_278 = 9'h116 == _GEN_7170 ? ram_278 : _GEN_277; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_279 = 9'h117 == _GEN_7170 ? ram_279 : _GEN_278; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_280 = 9'h118 == _GEN_7170 ? ram_280 : _GEN_279; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_281 = 9'h119 == _GEN_7170 ? ram_281 : _GEN_280; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_282 = 9'h11a == _GEN_7170 ? ram_282 : _GEN_281; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_283 = 9'h11b == _GEN_7170 ? ram_283 : _GEN_282; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_284 = 9'h11c == _GEN_7170 ? ram_284 : _GEN_283; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_285 = 9'h11d == _GEN_7170 ? ram_285 : _GEN_284; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_286 = 9'h11e == _GEN_7170 ? ram_286 : _GEN_285; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_287 = 9'h11f == _GEN_7170 ? ram_287 : _GEN_286; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_288 = 9'h120 == _GEN_7170 ? ram_288 : _GEN_287; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_289 = 9'h121 == _GEN_7170 ? ram_289 : _GEN_288; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_290 = 9'h122 == _GEN_7170 ? ram_290 : _GEN_289; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_291 = 9'h123 == _GEN_7170 ? ram_291 : _GEN_290; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_292 = 9'h124 == _GEN_7170 ? ram_292 : _GEN_291; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_293 = 9'h125 == _GEN_7170 ? ram_293 : _GEN_292; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_294 = 9'h126 == _GEN_7170 ? ram_294 : _GEN_293; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_295 = 9'h127 == _GEN_7170 ? ram_295 : _GEN_294; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_296 = 9'h128 == _GEN_7170 ? ram_296 : _GEN_295; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_297 = 9'h129 == _GEN_7170 ? ram_297 : _GEN_296; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_298 = 9'h12a == _GEN_7170 ? ram_298 : _GEN_297; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_299 = 9'h12b == _GEN_7170 ? ram_299 : _GEN_298; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_300 = 9'h12c == _GEN_7170 ? ram_300 : _GEN_299; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_301 = 9'h12d == _GEN_7170 ? ram_301 : _GEN_300; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_302 = 9'h12e == _GEN_7170 ? ram_302 : _GEN_301; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_303 = 9'h12f == _GEN_7170 ? ram_303 : _GEN_302; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_304 = 9'h130 == _GEN_7170 ? ram_304 : _GEN_303; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_305 = 9'h131 == _GEN_7170 ? ram_305 : _GEN_304; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_306 = 9'h132 == _GEN_7170 ? ram_306 : _GEN_305; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_307 = 9'h133 == _GEN_7170 ? ram_307 : _GEN_306; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_308 = 9'h134 == _GEN_7170 ? ram_308 : _GEN_307; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_309 = 9'h135 == _GEN_7170 ? ram_309 : _GEN_308; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_310 = 9'h136 == _GEN_7170 ? ram_310 : _GEN_309; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_311 = 9'h137 == _GEN_7170 ? ram_311 : _GEN_310; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_312 = 9'h138 == _GEN_7170 ? ram_312 : _GEN_311; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_313 = 9'h139 == _GEN_7170 ? ram_313 : _GEN_312; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_314 = 9'h13a == _GEN_7170 ? ram_314 : _GEN_313; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_315 = 9'h13b == _GEN_7170 ? ram_315 : _GEN_314; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_316 = 9'h13c == _GEN_7170 ? ram_316 : _GEN_315; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_317 = 9'h13d == _GEN_7170 ? ram_317 : _GEN_316; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_318 = 9'h13e == _GEN_7170 ? ram_318 : _GEN_317; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_319 = 9'h13f == _GEN_7170 ? ram_319 : _GEN_318; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_320 = 9'h140 == _GEN_7170 ? ram_320 : _GEN_319; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_321 = 9'h141 == _GEN_7170 ? ram_321 : _GEN_320; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_322 = 9'h142 == _GEN_7170 ? ram_322 : _GEN_321; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_323 = 9'h143 == _GEN_7170 ? ram_323 : _GEN_322; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_324 = 9'h144 == _GEN_7170 ? ram_324 : _GEN_323; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_325 = 9'h145 == _GEN_7170 ? ram_325 : _GEN_324; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_326 = 9'h146 == _GEN_7170 ? ram_326 : _GEN_325; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_327 = 9'h147 == _GEN_7170 ? ram_327 : _GEN_326; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_328 = 9'h148 == _GEN_7170 ? ram_328 : _GEN_327; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_329 = 9'h149 == _GEN_7170 ? ram_329 : _GEN_328; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_330 = 9'h14a == _GEN_7170 ? ram_330 : _GEN_329; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_331 = 9'h14b == _GEN_7170 ? ram_331 : _GEN_330; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_332 = 9'h14c == _GEN_7170 ? ram_332 : _GEN_331; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_333 = 9'h14d == _GEN_7170 ? ram_333 : _GEN_332; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_334 = 9'h14e == _GEN_7170 ? ram_334 : _GEN_333; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_335 = 9'h14f == _GEN_7170 ? ram_335 : _GEN_334; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_336 = 9'h150 == _GEN_7170 ? ram_336 : _GEN_335; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_337 = 9'h151 == _GEN_7170 ? ram_337 : _GEN_336; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_338 = 9'h152 == _GEN_7170 ? ram_338 : _GEN_337; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_339 = 9'h153 == _GEN_7170 ? ram_339 : _GEN_338; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_340 = 9'h154 == _GEN_7170 ? ram_340 : _GEN_339; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_341 = 9'h155 == _GEN_7170 ? ram_341 : _GEN_340; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_342 = 9'h156 == _GEN_7170 ? ram_342 : _GEN_341; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_343 = 9'h157 == _GEN_7170 ? ram_343 : _GEN_342; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_344 = 9'h158 == _GEN_7170 ? ram_344 : _GEN_343; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_345 = 9'h159 == _GEN_7170 ? ram_345 : _GEN_344; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_346 = 9'h15a == _GEN_7170 ? ram_346 : _GEN_345; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_347 = 9'h15b == _GEN_7170 ? ram_347 : _GEN_346; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_348 = 9'h15c == _GEN_7170 ? ram_348 : _GEN_347; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_349 = 9'h15d == _GEN_7170 ? ram_349 : _GEN_348; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_350 = 9'h15e == _GEN_7170 ? ram_350 : _GEN_349; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_351 = 9'h15f == _GEN_7170 ? ram_351 : _GEN_350; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_352 = 9'h160 == _GEN_7170 ? ram_352 : _GEN_351; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_353 = 9'h161 == _GEN_7170 ? ram_353 : _GEN_352; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_354 = 9'h162 == _GEN_7170 ? ram_354 : _GEN_353; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_355 = 9'h163 == _GEN_7170 ? ram_355 : _GEN_354; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_356 = 9'h164 == _GEN_7170 ? ram_356 : _GEN_355; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_357 = 9'h165 == _GEN_7170 ? ram_357 : _GEN_356; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_358 = 9'h166 == _GEN_7170 ? ram_358 : _GEN_357; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_359 = 9'h167 == _GEN_7170 ? ram_359 : _GEN_358; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_360 = 9'h168 == _GEN_7170 ? ram_360 : _GEN_359; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_361 = 9'h169 == _GEN_7170 ? ram_361 : _GEN_360; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_362 = 9'h16a == _GEN_7170 ? ram_362 : _GEN_361; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_363 = 9'h16b == _GEN_7170 ? ram_363 : _GEN_362; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_364 = 9'h16c == _GEN_7170 ? ram_364 : _GEN_363; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_365 = 9'h16d == _GEN_7170 ? ram_365 : _GEN_364; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_366 = 9'h16e == _GEN_7170 ? ram_366 : _GEN_365; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_367 = 9'h16f == _GEN_7170 ? ram_367 : _GEN_366; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_368 = 9'h170 == _GEN_7170 ? ram_368 : _GEN_367; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_369 = 9'h171 == _GEN_7170 ? ram_369 : _GEN_368; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_370 = 9'h172 == _GEN_7170 ? ram_370 : _GEN_369; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_371 = 9'h173 == _GEN_7170 ? ram_371 : _GEN_370; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_372 = 9'h174 == _GEN_7170 ? ram_372 : _GEN_371; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_373 = 9'h175 == _GEN_7170 ? ram_373 : _GEN_372; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_374 = 9'h176 == _GEN_7170 ? ram_374 : _GEN_373; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_375 = 9'h177 == _GEN_7170 ? ram_375 : _GEN_374; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_376 = 9'h178 == _GEN_7170 ? ram_376 : _GEN_375; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_377 = 9'h179 == _GEN_7170 ? ram_377 : _GEN_376; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_378 = 9'h17a == _GEN_7170 ? ram_378 : _GEN_377; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_379 = 9'h17b == _GEN_7170 ? ram_379 : _GEN_378; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_380 = 9'h17c == _GEN_7170 ? ram_380 : _GEN_379; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_381 = 9'h17d == _GEN_7170 ? ram_381 : _GEN_380; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_382 = 9'h17e == _GEN_7170 ? ram_382 : _GEN_381; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_383 = 9'h17f == _GEN_7170 ? ram_383 : _GEN_382; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_384 = 9'h180 == _GEN_7170 ? ram_384 : _GEN_383; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_385 = 9'h181 == _GEN_7170 ? ram_385 : _GEN_384; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_386 = 9'h182 == _GEN_7170 ? ram_386 : _GEN_385; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_387 = 9'h183 == _GEN_7170 ? ram_387 : _GEN_386; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_388 = 9'h184 == _GEN_7170 ? ram_388 : _GEN_387; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_389 = 9'h185 == _GEN_7170 ? ram_389 : _GEN_388; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_390 = 9'h186 == _GEN_7170 ? ram_390 : _GEN_389; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_391 = 9'h187 == _GEN_7170 ? ram_391 : _GEN_390; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_392 = 9'h188 == _GEN_7170 ? ram_392 : _GEN_391; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_393 = 9'h189 == _GEN_7170 ? ram_393 : _GEN_392; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_394 = 9'h18a == _GEN_7170 ? ram_394 : _GEN_393; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_395 = 9'h18b == _GEN_7170 ? ram_395 : _GEN_394; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_396 = 9'h18c == _GEN_7170 ? ram_396 : _GEN_395; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_397 = 9'h18d == _GEN_7170 ? ram_397 : _GEN_396; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_398 = 9'h18e == _GEN_7170 ? ram_398 : _GEN_397; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_399 = 9'h18f == _GEN_7170 ? ram_399 : _GEN_398; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_400 = 9'h190 == _GEN_7170 ? ram_400 : _GEN_399; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_401 = 9'h191 == _GEN_7170 ? ram_401 : _GEN_400; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_402 = 9'h192 == _GEN_7170 ? ram_402 : _GEN_401; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_403 = 9'h193 == _GEN_7170 ? ram_403 : _GEN_402; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_404 = 9'h194 == _GEN_7170 ? ram_404 : _GEN_403; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_405 = 9'h195 == _GEN_7170 ? ram_405 : _GEN_404; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_406 = 9'h196 == _GEN_7170 ? ram_406 : _GEN_405; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_407 = 9'h197 == _GEN_7170 ? ram_407 : _GEN_406; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_408 = 9'h198 == _GEN_7170 ? ram_408 : _GEN_407; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_409 = 9'h199 == _GEN_7170 ? ram_409 : _GEN_408; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_410 = 9'h19a == _GEN_7170 ? ram_410 : _GEN_409; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_411 = 9'h19b == _GEN_7170 ? ram_411 : _GEN_410; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_412 = 9'h19c == _GEN_7170 ? ram_412 : _GEN_411; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_413 = 9'h19d == _GEN_7170 ? ram_413 : _GEN_412; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_414 = 9'h19e == _GEN_7170 ? ram_414 : _GEN_413; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_415 = 9'h19f == _GEN_7170 ? ram_415 : _GEN_414; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_416 = 9'h1a0 == _GEN_7170 ? ram_416 : _GEN_415; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_417 = 9'h1a1 == _GEN_7170 ? ram_417 : _GEN_416; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_418 = 9'h1a2 == _GEN_7170 ? ram_418 : _GEN_417; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_419 = 9'h1a3 == _GEN_7170 ? ram_419 : _GEN_418; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_420 = 9'h1a4 == _GEN_7170 ? ram_420 : _GEN_419; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_421 = 9'h1a5 == _GEN_7170 ? ram_421 : _GEN_420; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_422 = 9'h1a6 == _GEN_7170 ? ram_422 : _GEN_421; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_423 = 9'h1a7 == _GEN_7170 ? ram_423 : _GEN_422; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_424 = 9'h1a8 == _GEN_7170 ? ram_424 : _GEN_423; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_425 = 9'h1a9 == _GEN_7170 ? ram_425 : _GEN_424; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_426 = 9'h1aa == _GEN_7170 ? ram_426 : _GEN_425; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_427 = 9'h1ab == _GEN_7170 ? ram_427 : _GEN_426; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_428 = 9'h1ac == _GEN_7170 ? ram_428 : _GEN_427; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_429 = 9'h1ad == _GEN_7170 ? ram_429 : _GEN_428; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_430 = 9'h1ae == _GEN_7170 ? ram_430 : _GEN_429; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_431 = 9'h1af == _GEN_7170 ? ram_431 : _GEN_430; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_432 = 9'h1b0 == _GEN_7170 ? ram_432 : _GEN_431; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_433 = 9'h1b1 == _GEN_7170 ? ram_433 : _GEN_432; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_434 = 9'h1b2 == _GEN_7170 ? ram_434 : _GEN_433; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_435 = 9'h1b3 == _GEN_7170 ? ram_435 : _GEN_434; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_436 = 9'h1b4 == _GEN_7170 ? ram_436 : _GEN_435; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_437 = 9'h1b5 == _GEN_7170 ? ram_437 : _GEN_436; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_438 = 9'h1b6 == _GEN_7170 ? ram_438 : _GEN_437; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_439 = 9'h1b7 == _GEN_7170 ? ram_439 : _GEN_438; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_440 = 9'h1b8 == _GEN_7170 ? ram_440 : _GEN_439; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_441 = 9'h1b9 == _GEN_7170 ? ram_441 : _GEN_440; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_442 = 9'h1ba == _GEN_7170 ? ram_442 : _GEN_441; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_443 = 9'h1bb == _GEN_7170 ? ram_443 : _GEN_442; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_444 = 9'h1bc == _GEN_7170 ? ram_444 : _GEN_443; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_445 = 9'h1bd == _GEN_7170 ? ram_445 : _GEN_444; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_446 = 9'h1be == _GEN_7170 ? ram_446 : _GEN_445; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_447 = 9'h1bf == _GEN_7170 ? ram_447 : _GEN_446; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_448 = 9'h1c0 == _GEN_7170 ? ram_448 : _GEN_447; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_449 = 9'h1c1 == _GEN_7170 ? ram_449 : _GEN_448; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_450 = 9'h1c2 == _GEN_7170 ? ram_450 : _GEN_449; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_451 = 9'h1c3 == _GEN_7170 ? ram_451 : _GEN_450; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_452 = 9'h1c4 == _GEN_7170 ? ram_452 : _GEN_451; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_453 = 9'h1c5 == _GEN_7170 ? ram_453 : _GEN_452; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_454 = 9'h1c6 == _GEN_7170 ? ram_454 : _GEN_453; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_455 = 9'h1c7 == _GEN_7170 ? ram_455 : _GEN_454; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_456 = 9'h1c8 == _GEN_7170 ? ram_456 : _GEN_455; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_457 = 9'h1c9 == _GEN_7170 ? ram_457 : _GEN_456; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_458 = 9'h1ca == _GEN_7170 ? ram_458 : _GEN_457; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_459 = 9'h1cb == _GEN_7170 ? ram_459 : _GEN_458; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_460 = 9'h1cc == _GEN_7170 ? ram_460 : _GEN_459; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_461 = 9'h1cd == _GEN_7170 ? ram_461 : _GEN_460; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_462 = 9'h1ce == _GEN_7170 ? ram_462 : _GEN_461; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_463 = 9'h1cf == _GEN_7170 ? ram_463 : _GEN_462; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_464 = 9'h1d0 == _GEN_7170 ? ram_464 : _GEN_463; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_465 = 9'h1d1 == _GEN_7170 ? ram_465 : _GEN_464; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_466 = 9'h1d2 == _GEN_7170 ? ram_466 : _GEN_465; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_467 = 9'h1d3 == _GEN_7170 ? ram_467 : _GEN_466; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_468 = 9'h1d4 == _GEN_7170 ? ram_468 : _GEN_467; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_469 = 9'h1d5 == _GEN_7170 ? ram_469 : _GEN_468; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_470 = 9'h1d6 == _GEN_7170 ? ram_470 : _GEN_469; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_471 = 9'h1d7 == _GEN_7170 ? ram_471 : _GEN_470; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_472 = 9'h1d8 == _GEN_7170 ? ram_472 : _GEN_471; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_473 = 9'h1d9 == _GEN_7170 ? ram_473 : _GEN_472; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_474 = 9'h1da == _GEN_7170 ? ram_474 : _GEN_473; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_475 = 9'h1db == _GEN_7170 ? ram_475 : _GEN_474; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_476 = 9'h1dc == _GEN_7170 ? ram_476 : _GEN_475; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_477 = 9'h1dd == _GEN_7170 ? ram_477 : _GEN_476; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_478 = 9'h1de == _GEN_7170 ? ram_478 : _GEN_477; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_479 = 9'h1df == _GEN_7170 ? ram_479 : _GEN_478; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_480 = 9'h1e0 == _GEN_7170 ? ram_480 : _GEN_479; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_481 = 9'h1e1 == _GEN_7170 ? ram_481 : _GEN_480; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_482 = 9'h1e2 == _GEN_7170 ? ram_482 : _GEN_481; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_483 = 9'h1e3 == _GEN_7170 ? ram_483 : _GEN_482; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_484 = 9'h1e4 == _GEN_7170 ? ram_484 : _GEN_483; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_485 = 9'h1e5 == _GEN_7170 ? ram_485 : _GEN_484; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_486 = 9'h1e6 == _GEN_7170 ? ram_486 : _GEN_485; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_487 = 9'h1e7 == _GEN_7170 ? ram_487 : _GEN_486; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_488 = 9'h1e8 == _GEN_7170 ? ram_488 : _GEN_487; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_489 = 9'h1e9 == _GEN_7170 ? ram_489 : _GEN_488; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_490 = 9'h1ea == _GEN_7170 ? ram_490 : _GEN_489; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_491 = 9'h1eb == _GEN_7170 ? ram_491 : _GEN_490; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_492 = 9'h1ec == _GEN_7170 ? ram_492 : _GEN_491; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_493 = 9'h1ed == _GEN_7170 ? ram_493 : _GEN_492; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_494 = 9'h1ee == _GEN_7170 ? ram_494 : _GEN_493; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_495 = 9'h1ef == _GEN_7170 ? ram_495 : _GEN_494; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_496 = 9'h1f0 == _GEN_7170 ? ram_496 : _GEN_495; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_497 = 9'h1f1 == _GEN_7170 ? ram_497 : _GEN_496; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_498 = 9'h1f2 == _GEN_7170 ? ram_498 : _GEN_497; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_499 = 9'h1f3 == _GEN_7170 ? ram_499 : _GEN_498; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_500 = 9'h1f4 == _GEN_7170 ? ram_500 : _GEN_499; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_501 = 9'h1f5 == _GEN_7170 ? ram_501 : _GEN_500; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_502 = 9'h1f6 == _GEN_7170 ? ram_502 : _GEN_501; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_503 = 9'h1f7 == _GEN_7170 ? ram_503 : _GEN_502; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_504 = 9'h1f8 == _GEN_7170 ? ram_504 : _GEN_503; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_505 = 9'h1f9 == _GEN_7170 ? ram_505 : _GEN_504; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_506 = 9'h1fa == _GEN_7170 ? ram_506 : _GEN_505; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_507 = 9'h1fb == _GEN_7170 ? ram_507 : _GEN_506; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_508 = 9'h1fc == _GEN_7170 ? ram_508 : _GEN_507; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_509 = 9'h1fd == _GEN_7170 ? ram_509 : _GEN_508; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_510 = 9'h1fe == _GEN_7170 ? ram_510 : _GEN_509; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_511 = 9'h1ff == _GEN_7170 ? ram_511 : _GEN_510; // @[DataMemory.scala 42:{28,28}]
  wire [9:0] _GEN_7426 = {{2'd0}, io_addr[9:2]}; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_512 = 10'h200 == _GEN_7426 ? ram_512 : _GEN_511; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_513 = 10'h201 == _GEN_7426 ? ram_513 : _GEN_512; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_514 = 10'h202 == _GEN_7426 ? ram_514 : _GEN_513; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_515 = 10'h203 == _GEN_7426 ? ram_515 : _GEN_514; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_516 = 10'h204 == _GEN_7426 ? ram_516 : _GEN_515; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_517 = 10'h205 == _GEN_7426 ? ram_517 : _GEN_516; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_518 = 10'h206 == _GEN_7426 ? ram_518 : _GEN_517; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_519 = 10'h207 == _GEN_7426 ? ram_519 : _GEN_518; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_520 = 10'h208 == _GEN_7426 ? ram_520 : _GEN_519; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_521 = 10'h209 == _GEN_7426 ? ram_521 : _GEN_520; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_522 = 10'h20a == _GEN_7426 ? ram_522 : _GEN_521; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_523 = 10'h20b == _GEN_7426 ? ram_523 : _GEN_522; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_524 = 10'h20c == _GEN_7426 ? ram_524 : _GEN_523; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_525 = 10'h20d == _GEN_7426 ? ram_525 : _GEN_524; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_526 = 10'h20e == _GEN_7426 ? ram_526 : _GEN_525; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_527 = 10'h20f == _GEN_7426 ? ram_527 : _GEN_526; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_528 = 10'h210 == _GEN_7426 ? ram_528 : _GEN_527; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_529 = 10'h211 == _GEN_7426 ? ram_529 : _GEN_528; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_530 = 10'h212 == _GEN_7426 ? ram_530 : _GEN_529; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_531 = 10'h213 == _GEN_7426 ? ram_531 : _GEN_530; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_532 = 10'h214 == _GEN_7426 ? ram_532 : _GEN_531; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_533 = 10'h215 == _GEN_7426 ? ram_533 : _GEN_532; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_534 = 10'h216 == _GEN_7426 ? ram_534 : _GEN_533; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_535 = 10'h217 == _GEN_7426 ? ram_535 : _GEN_534; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_536 = 10'h218 == _GEN_7426 ? ram_536 : _GEN_535; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_537 = 10'h219 == _GEN_7426 ? ram_537 : _GEN_536; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_538 = 10'h21a == _GEN_7426 ? ram_538 : _GEN_537; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_539 = 10'h21b == _GEN_7426 ? ram_539 : _GEN_538; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_540 = 10'h21c == _GEN_7426 ? ram_540 : _GEN_539; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_541 = 10'h21d == _GEN_7426 ? ram_541 : _GEN_540; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_542 = 10'h21e == _GEN_7426 ? ram_542 : _GEN_541; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_543 = 10'h21f == _GEN_7426 ? ram_543 : _GEN_542; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_544 = 10'h220 == _GEN_7426 ? ram_544 : _GEN_543; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_545 = 10'h221 == _GEN_7426 ? ram_545 : _GEN_544; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_546 = 10'h222 == _GEN_7426 ? ram_546 : _GEN_545; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_547 = 10'h223 == _GEN_7426 ? ram_547 : _GEN_546; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_548 = 10'h224 == _GEN_7426 ? ram_548 : _GEN_547; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_549 = 10'h225 == _GEN_7426 ? ram_549 : _GEN_548; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_550 = 10'h226 == _GEN_7426 ? ram_550 : _GEN_549; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_551 = 10'h227 == _GEN_7426 ? ram_551 : _GEN_550; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_552 = 10'h228 == _GEN_7426 ? ram_552 : _GEN_551; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_553 = 10'h229 == _GEN_7426 ? ram_553 : _GEN_552; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_554 = 10'h22a == _GEN_7426 ? ram_554 : _GEN_553; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_555 = 10'h22b == _GEN_7426 ? ram_555 : _GEN_554; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_556 = 10'h22c == _GEN_7426 ? ram_556 : _GEN_555; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_557 = 10'h22d == _GEN_7426 ? ram_557 : _GEN_556; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_558 = 10'h22e == _GEN_7426 ? ram_558 : _GEN_557; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_559 = 10'h22f == _GEN_7426 ? ram_559 : _GEN_558; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_560 = 10'h230 == _GEN_7426 ? ram_560 : _GEN_559; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_561 = 10'h231 == _GEN_7426 ? ram_561 : _GEN_560; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_562 = 10'h232 == _GEN_7426 ? ram_562 : _GEN_561; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_563 = 10'h233 == _GEN_7426 ? ram_563 : _GEN_562; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_564 = 10'h234 == _GEN_7426 ? ram_564 : _GEN_563; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_565 = 10'h235 == _GEN_7426 ? ram_565 : _GEN_564; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_566 = 10'h236 == _GEN_7426 ? ram_566 : _GEN_565; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_567 = 10'h237 == _GEN_7426 ? ram_567 : _GEN_566; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_568 = 10'h238 == _GEN_7426 ? ram_568 : _GEN_567; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_569 = 10'h239 == _GEN_7426 ? ram_569 : _GEN_568; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_570 = 10'h23a == _GEN_7426 ? ram_570 : _GEN_569; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_571 = 10'h23b == _GEN_7426 ? ram_571 : _GEN_570; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_572 = 10'h23c == _GEN_7426 ? ram_572 : _GEN_571; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_573 = 10'h23d == _GEN_7426 ? ram_573 : _GEN_572; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_574 = 10'h23e == _GEN_7426 ? ram_574 : _GEN_573; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_575 = 10'h23f == _GEN_7426 ? ram_575 : _GEN_574; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_576 = 10'h240 == _GEN_7426 ? ram_576 : _GEN_575; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_577 = 10'h241 == _GEN_7426 ? ram_577 : _GEN_576; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_578 = 10'h242 == _GEN_7426 ? ram_578 : _GEN_577; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_579 = 10'h243 == _GEN_7426 ? ram_579 : _GEN_578; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_580 = 10'h244 == _GEN_7426 ? ram_580 : _GEN_579; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_581 = 10'h245 == _GEN_7426 ? ram_581 : _GEN_580; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_582 = 10'h246 == _GEN_7426 ? ram_582 : _GEN_581; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_583 = 10'h247 == _GEN_7426 ? ram_583 : _GEN_582; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_584 = 10'h248 == _GEN_7426 ? ram_584 : _GEN_583; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_585 = 10'h249 == _GEN_7426 ? ram_585 : _GEN_584; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_586 = 10'h24a == _GEN_7426 ? ram_586 : _GEN_585; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_587 = 10'h24b == _GEN_7426 ? ram_587 : _GEN_586; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_588 = 10'h24c == _GEN_7426 ? ram_588 : _GEN_587; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_589 = 10'h24d == _GEN_7426 ? ram_589 : _GEN_588; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_590 = 10'h24e == _GEN_7426 ? ram_590 : _GEN_589; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_591 = 10'h24f == _GEN_7426 ? ram_591 : _GEN_590; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_592 = 10'h250 == _GEN_7426 ? ram_592 : _GEN_591; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_593 = 10'h251 == _GEN_7426 ? ram_593 : _GEN_592; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_594 = 10'h252 == _GEN_7426 ? ram_594 : _GEN_593; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_595 = 10'h253 == _GEN_7426 ? ram_595 : _GEN_594; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_596 = 10'h254 == _GEN_7426 ? ram_596 : _GEN_595; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_597 = 10'h255 == _GEN_7426 ? ram_597 : _GEN_596; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_598 = 10'h256 == _GEN_7426 ? ram_598 : _GEN_597; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_599 = 10'h257 == _GEN_7426 ? ram_599 : _GEN_598; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_600 = 10'h258 == _GEN_7426 ? ram_600 : _GEN_599; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_601 = 10'h259 == _GEN_7426 ? ram_601 : _GEN_600; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_602 = 10'h25a == _GEN_7426 ? ram_602 : _GEN_601; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_603 = 10'h25b == _GEN_7426 ? ram_603 : _GEN_602; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_604 = 10'h25c == _GEN_7426 ? ram_604 : _GEN_603; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_605 = 10'h25d == _GEN_7426 ? ram_605 : _GEN_604; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_606 = 10'h25e == _GEN_7426 ? ram_606 : _GEN_605; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_607 = 10'h25f == _GEN_7426 ? ram_607 : _GEN_606; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_608 = 10'h260 == _GEN_7426 ? ram_608 : _GEN_607; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_609 = 10'h261 == _GEN_7426 ? ram_609 : _GEN_608; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_610 = 10'h262 == _GEN_7426 ? ram_610 : _GEN_609; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_611 = 10'h263 == _GEN_7426 ? ram_611 : _GEN_610; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_612 = 10'h264 == _GEN_7426 ? ram_612 : _GEN_611; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_613 = 10'h265 == _GEN_7426 ? ram_613 : _GEN_612; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_614 = 10'h266 == _GEN_7426 ? ram_614 : _GEN_613; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_615 = 10'h267 == _GEN_7426 ? ram_615 : _GEN_614; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_616 = 10'h268 == _GEN_7426 ? ram_616 : _GEN_615; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_617 = 10'h269 == _GEN_7426 ? ram_617 : _GEN_616; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_618 = 10'h26a == _GEN_7426 ? ram_618 : _GEN_617; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_619 = 10'h26b == _GEN_7426 ? ram_619 : _GEN_618; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_620 = 10'h26c == _GEN_7426 ? ram_620 : _GEN_619; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_621 = 10'h26d == _GEN_7426 ? ram_621 : _GEN_620; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_622 = 10'h26e == _GEN_7426 ? ram_622 : _GEN_621; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_623 = 10'h26f == _GEN_7426 ? ram_623 : _GEN_622; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_624 = 10'h270 == _GEN_7426 ? ram_624 : _GEN_623; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_625 = 10'h271 == _GEN_7426 ? ram_625 : _GEN_624; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_626 = 10'h272 == _GEN_7426 ? ram_626 : _GEN_625; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_627 = 10'h273 == _GEN_7426 ? ram_627 : _GEN_626; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_628 = 10'h274 == _GEN_7426 ? ram_628 : _GEN_627; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_629 = 10'h275 == _GEN_7426 ? ram_629 : _GEN_628; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_630 = 10'h276 == _GEN_7426 ? ram_630 : _GEN_629; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_631 = 10'h277 == _GEN_7426 ? ram_631 : _GEN_630; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_632 = 10'h278 == _GEN_7426 ? ram_632 : _GEN_631; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_633 = 10'h279 == _GEN_7426 ? ram_633 : _GEN_632; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_634 = 10'h27a == _GEN_7426 ? ram_634 : _GEN_633; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_635 = 10'h27b == _GEN_7426 ? ram_635 : _GEN_634; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_636 = 10'h27c == _GEN_7426 ? ram_636 : _GEN_635; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_637 = 10'h27d == _GEN_7426 ? ram_637 : _GEN_636; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_638 = 10'h27e == _GEN_7426 ? ram_638 : _GEN_637; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_639 = 10'h27f == _GEN_7426 ? ram_639 : _GEN_638; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_640 = 10'h280 == _GEN_7426 ? ram_640 : _GEN_639; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_641 = 10'h281 == _GEN_7426 ? ram_641 : _GEN_640; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_642 = 10'h282 == _GEN_7426 ? ram_642 : _GEN_641; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_643 = 10'h283 == _GEN_7426 ? ram_643 : _GEN_642; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_644 = 10'h284 == _GEN_7426 ? ram_644 : _GEN_643; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_645 = 10'h285 == _GEN_7426 ? ram_645 : _GEN_644; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_646 = 10'h286 == _GEN_7426 ? ram_646 : _GEN_645; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_647 = 10'h287 == _GEN_7426 ? ram_647 : _GEN_646; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_648 = 10'h288 == _GEN_7426 ? ram_648 : _GEN_647; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_649 = 10'h289 == _GEN_7426 ? ram_649 : _GEN_648; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_650 = 10'h28a == _GEN_7426 ? ram_650 : _GEN_649; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_651 = 10'h28b == _GEN_7426 ? ram_651 : _GEN_650; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_652 = 10'h28c == _GEN_7426 ? ram_652 : _GEN_651; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_653 = 10'h28d == _GEN_7426 ? ram_653 : _GEN_652; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_654 = 10'h28e == _GEN_7426 ? ram_654 : _GEN_653; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_655 = 10'h28f == _GEN_7426 ? ram_655 : _GEN_654; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_656 = 10'h290 == _GEN_7426 ? ram_656 : _GEN_655; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_657 = 10'h291 == _GEN_7426 ? ram_657 : _GEN_656; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_658 = 10'h292 == _GEN_7426 ? ram_658 : _GEN_657; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_659 = 10'h293 == _GEN_7426 ? ram_659 : _GEN_658; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_660 = 10'h294 == _GEN_7426 ? ram_660 : _GEN_659; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_661 = 10'h295 == _GEN_7426 ? ram_661 : _GEN_660; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_662 = 10'h296 == _GEN_7426 ? ram_662 : _GEN_661; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_663 = 10'h297 == _GEN_7426 ? ram_663 : _GEN_662; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_664 = 10'h298 == _GEN_7426 ? ram_664 : _GEN_663; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_665 = 10'h299 == _GEN_7426 ? ram_665 : _GEN_664; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_666 = 10'h29a == _GEN_7426 ? ram_666 : _GEN_665; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_667 = 10'h29b == _GEN_7426 ? ram_667 : _GEN_666; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_668 = 10'h29c == _GEN_7426 ? ram_668 : _GEN_667; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_669 = 10'h29d == _GEN_7426 ? ram_669 : _GEN_668; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_670 = 10'h29e == _GEN_7426 ? ram_670 : _GEN_669; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_671 = 10'h29f == _GEN_7426 ? ram_671 : _GEN_670; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_672 = 10'h2a0 == _GEN_7426 ? ram_672 : _GEN_671; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_673 = 10'h2a1 == _GEN_7426 ? ram_673 : _GEN_672; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_674 = 10'h2a2 == _GEN_7426 ? ram_674 : _GEN_673; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_675 = 10'h2a3 == _GEN_7426 ? ram_675 : _GEN_674; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_676 = 10'h2a4 == _GEN_7426 ? ram_676 : _GEN_675; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_677 = 10'h2a5 == _GEN_7426 ? ram_677 : _GEN_676; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_678 = 10'h2a6 == _GEN_7426 ? ram_678 : _GEN_677; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_679 = 10'h2a7 == _GEN_7426 ? ram_679 : _GEN_678; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_680 = 10'h2a8 == _GEN_7426 ? ram_680 : _GEN_679; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_681 = 10'h2a9 == _GEN_7426 ? ram_681 : _GEN_680; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_682 = 10'h2aa == _GEN_7426 ? ram_682 : _GEN_681; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_683 = 10'h2ab == _GEN_7426 ? ram_683 : _GEN_682; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_684 = 10'h2ac == _GEN_7426 ? ram_684 : _GEN_683; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_685 = 10'h2ad == _GEN_7426 ? ram_685 : _GEN_684; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_686 = 10'h2ae == _GEN_7426 ? ram_686 : _GEN_685; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_687 = 10'h2af == _GEN_7426 ? ram_687 : _GEN_686; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_688 = 10'h2b0 == _GEN_7426 ? ram_688 : _GEN_687; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_689 = 10'h2b1 == _GEN_7426 ? ram_689 : _GEN_688; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_690 = 10'h2b2 == _GEN_7426 ? ram_690 : _GEN_689; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_691 = 10'h2b3 == _GEN_7426 ? ram_691 : _GEN_690; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_692 = 10'h2b4 == _GEN_7426 ? ram_692 : _GEN_691; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_693 = 10'h2b5 == _GEN_7426 ? ram_693 : _GEN_692; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_694 = 10'h2b6 == _GEN_7426 ? ram_694 : _GEN_693; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_695 = 10'h2b7 == _GEN_7426 ? ram_695 : _GEN_694; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_696 = 10'h2b8 == _GEN_7426 ? ram_696 : _GEN_695; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_697 = 10'h2b9 == _GEN_7426 ? ram_697 : _GEN_696; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_698 = 10'h2ba == _GEN_7426 ? ram_698 : _GEN_697; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_699 = 10'h2bb == _GEN_7426 ? ram_699 : _GEN_698; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_700 = 10'h2bc == _GEN_7426 ? ram_700 : _GEN_699; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_701 = 10'h2bd == _GEN_7426 ? ram_701 : _GEN_700; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_702 = 10'h2be == _GEN_7426 ? ram_702 : _GEN_701; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_703 = 10'h2bf == _GEN_7426 ? ram_703 : _GEN_702; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_704 = 10'h2c0 == _GEN_7426 ? ram_704 : _GEN_703; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_705 = 10'h2c1 == _GEN_7426 ? ram_705 : _GEN_704; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_706 = 10'h2c2 == _GEN_7426 ? ram_706 : _GEN_705; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_707 = 10'h2c3 == _GEN_7426 ? ram_707 : _GEN_706; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_708 = 10'h2c4 == _GEN_7426 ? ram_708 : _GEN_707; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_709 = 10'h2c5 == _GEN_7426 ? ram_709 : _GEN_708; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_710 = 10'h2c6 == _GEN_7426 ? ram_710 : _GEN_709; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_711 = 10'h2c7 == _GEN_7426 ? ram_711 : _GEN_710; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_712 = 10'h2c8 == _GEN_7426 ? ram_712 : _GEN_711; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_713 = 10'h2c9 == _GEN_7426 ? ram_713 : _GEN_712; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_714 = 10'h2ca == _GEN_7426 ? ram_714 : _GEN_713; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_715 = 10'h2cb == _GEN_7426 ? ram_715 : _GEN_714; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_716 = 10'h2cc == _GEN_7426 ? ram_716 : _GEN_715; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_717 = 10'h2cd == _GEN_7426 ? ram_717 : _GEN_716; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_718 = 10'h2ce == _GEN_7426 ? ram_718 : _GEN_717; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_719 = 10'h2cf == _GEN_7426 ? ram_719 : _GEN_718; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_720 = 10'h2d0 == _GEN_7426 ? ram_720 : _GEN_719; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_721 = 10'h2d1 == _GEN_7426 ? ram_721 : _GEN_720; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_722 = 10'h2d2 == _GEN_7426 ? ram_722 : _GEN_721; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_723 = 10'h2d3 == _GEN_7426 ? ram_723 : _GEN_722; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_724 = 10'h2d4 == _GEN_7426 ? ram_724 : _GEN_723; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_725 = 10'h2d5 == _GEN_7426 ? ram_725 : _GEN_724; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_726 = 10'h2d6 == _GEN_7426 ? ram_726 : _GEN_725; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_727 = 10'h2d7 == _GEN_7426 ? ram_727 : _GEN_726; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_728 = 10'h2d8 == _GEN_7426 ? ram_728 : _GEN_727; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_729 = 10'h2d9 == _GEN_7426 ? ram_729 : _GEN_728; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_730 = 10'h2da == _GEN_7426 ? ram_730 : _GEN_729; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_731 = 10'h2db == _GEN_7426 ? ram_731 : _GEN_730; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_732 = 10'h2dc == _GEN_7426 ? ram_732 : _GEN_731; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_733 = 10'h2dd == _GEN_7426 ? ram_733 : _GEN_732; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_734 = 10'h2de == _GEN_7426 ? ram_734 : _GEN_733; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_735 = 10'h2df == _GEN_7426 ? ram_735 : _GEN_734; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_736 = 10'h2e0 == _GEN_7426 ? ram_736 : _GEN_735; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_737 = 10'h2e1 == _GEN_7426 ? ram_737 : _GEN_736; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_738 = 10'h2e2 == _GEN_7426 ? ram_738 : _GEN_737; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_739 = 10'h2e3 == _GEN_7426 ? ram_739 : _GEN_738; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_740 = 10'h2e4 == _GEN_7426 ? ram_740 : _GEN_739; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_741 = 10'h2e5 == _GEN_7426 ? ram_741 : _GEN_740; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_742 = 10'h2e6 == _GEN_7426 ? ram_742 : _GEN_741; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_743 = 10'h2e7 == _GEN_7426 ? ram_743 : _GEN_742; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_744 = 10'h2e8 == _GEN_7426 ? ram_744 : _GEN_743; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_745 = 10'h2e9 == _GEN_7426 ? ram_745 : _GEN_744; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_746 = 10'h2ea == _GEN_7426 ? ram_746 : _GEN_745; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_747 = 10'h2eb == _GEN_7426 ? ram_747 : _GEN_746; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_748 = 10'h2ec == _GEN_7426 ? ram_748 : _GEN_747; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_749 = 10'h2ed == _GEN_7426 ? ram_749 : _GEN_748; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_750 = 10'h2ee == _GEN_7426 ? ram_750 : _GEN_749; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_751 = 10'h2ef == _GEN_7426 ? ram_751 : _GEN_750; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_752 = 10'h2f0 == _GEN_7426 ? ram_752 : _GEN_751; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_753 = 10'h2f1 == _GEN_7426 ? ram_753 : _GEN_752; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_754 = 10'h2f2 == _GEN_7426 ? ram_754 : _GEN_753; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_755 = 10'h2f3 == _GEN_7426 ? ram_755 : _GEN_754; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_756 = 10'h2f4 == _GEN_7426 ? ram_756 : _GEN_755; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_757 = 10'h2f5 == _GEN_7426 ? ram_757 : _GEN_756; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_758 = 10'h2f6 == _GEN_7426 ? ram_758 : _GEN_757; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_759 = 10'h2f7 == _GEN_7426 ? ram_759 : _GEN_758; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_760 = 10'h2f8 == _GEN_7426 ? ram_760 : _GEN_759; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_761 = 10'h2f9 == _GEN_7426 ? ram_761 : _GEN_760; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_762 = 10'h2fa == _GEN_7426 ? ram_762 : _GEN_761; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_763 = 10'h2fb == _GEN_7426 ? ram_763 : _GEN_762; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_764 = 10'h2fc == _GEN_7426 ? ram_764 : _GEN_763; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_765 = 10'h2fd == _GEN_7426 ? ram_765 : _GEN_764; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_766 = 10'h2fe == _GEN_7426 ? ram_766 : _GEN_765; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_767 = 10'h2ff == _GEN_7426 ? ram_767 : _GEN_766; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_768 = 10'h300 == _GEN_7426 ? ram_768 : _GEN_767; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_769 = 10'h301 == _GEN_7426 ? ram_769 : _GEN_768; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_770 = 10'h302 == _GEN_7426 ? ram_770 : _GEN_769; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_771 = 10'h303 == _GEN_7426 ? ram_771 : _GEN_770; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_772 = 10'h304 == _GEN_7426 ? ram_772 : _GEN_771; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_773 = 10'h305 == _GEN_7426 ? ram_773 : _GEN_772; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_774 = 10'h306 == _GEN_7426 ? ram_774 : _GEN_773; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_775 = 10'h307 == _GEN_7426 ? ram_775 : _GEN_774; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_776 = 10'h308 == _GEN_7426 ? ram_776 : _GEN_775; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_777 = 10'h309 == _GEN_7426 ? ram_777 : _GEN_776; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_778 = 10'h30a == _GEN_7426 ? ram_778 : _GEN_777; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_779 = 10'h30b == _GEN_7426 ? ram_779 : _GEN_778; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_780 = 10'h30c == _GEN_7426 ? ram_780 : _GEN_779; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_781 = 10'h30d == _GEN_7426 ? ram_781 : _GEN_780; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_782 = 10'h30e == _GEN_7426 ? ram_782 : _GEN_781; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_783 = 10'h30f == _GEN_7426 ? ram_783 : _GEN_782; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_784 = 10'h310 == _GEN_7426 ? ram_784 : _GEN_783; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_785 = 10'h311 == _GEN_7426 ? ram_785 : _GEN_784; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_786 = 10'h312 == _GEN_7426 ? ram_786 : _GEN_785; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_787 = 10'h313 == _GEN_7426 ? ram_787 : _GEN_786; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_788 = 10'h314 == _GEN_7426 ? ram_788 : _GEN_787; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_789 = 10'h315 == _GEN_7426 ? ram_789 : _GEN_788; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_790 = 10'h316 == _GEN_7426 ? ram_790 : _GEN_789; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_791 = 10'h317 == _GEN_7426 ? ram_791 : _GEN_790; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_792 = 10'h318 == _GEN_7426 ? ram_792 : _GEN_791; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_793 = 10'h319 == _GEN_7426 ? ram_793 : _GEN_792; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_794 = 10'h31a == _GEN_7426 ? ram_794 : _GEN_793; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_795 = 10'h31b == _GEN_7426 ? ram_795 : _GEN_794; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_796 = 10'h31c == _GEN_7426 ? ram_796 : _GEN_795; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_797 = 10'h31d == _GEN_7426 ? ram_797 : _GEN_796; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_798 = 10'h31e == _GEN_7426 ? ram_798 : _GEN_797; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_799 = 10'h31f == _GEN_7426 ? ram_799 : _GEN_798; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_800 = 10'h320 == _GEN_7426 ? ram_800 : _GEN_799; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_801 = 10'h321 == _GEN_7426 ? ram_801 : _GEN_800; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_802 = 10'h322 == _GEN_7426 ? ram_802 : _GEN_801; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_803 = 10'h323 == _GEN_7426 ? ram_803 : _GEN_802; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_804 = 10'h324 == _GEN_7426 ? ram_804 : _GEN_803; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_805 = 10'h325 == _GEN_7426 ? ram_805 : _GEN_804; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_806 = 10'h326 == _GEN_7426 ? ram_806 : _GEN_805; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_807 = 10'h327 == _GEN_7426 ? ram_807 : _GEN_806; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_808 = 10'h328 == _GEN_7426 ? ram_808 : _GEN_807; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_809 = 10'h329 == _GEN_7426 ? ram_809 : _GEN_808; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_810 = 10'h32a == _GEN_7426 ? ram_810 : _GEN_809; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_811 = 10'h32b == _GEN_7426 ? ram_811 : _GEN_810; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_812 = 10'h32c == _GEN_7426 ? ram_812 : _GEN_811; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_813 = 10'h32d == _GEN_7426 ? ram_813 : _GEN_812; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_814 = 10'h32e == _GEN_7426 ? ram_814 : _GEN_813; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_815 = 10'h32f == _GEN_7426 ? ram_815 : _GEN_814; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_816 = 10'h330 == _GEN_7426 ? ram_816 : _GEN_815; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_817 = 10'h331 == _GEN_7426 ? ram_817 : _GEN_816; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_818 = 10'h332 == _GEN_7426 ? ram_818 : _GEN_817; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_819 = 10'h333 == _GEN_7426 ? ram_819 : _GEN_818; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_820 = 10'h334 == _GEN_7426 ? ram_820 : _GEN_819; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_821 = 10'h335 == _GEN_7426 ? ram_821 : _GEN_820; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_822 = 10'h336 == _GEN_7426 ? ram_822 : _GEN_821; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_823 = 10'h337 == _GEN_7426 ? ram_823 : _GEN_822; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_824 = 10'h338 == _GEN_7426 ? ram_824 : _GEN_823; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_825 = 10'h339 == _GEN_7426 ? ram_825 : _GEN_824; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_826 = 10'h33a == _GEN_7426 ? ram_826 : _GEN_825; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_827 = 10'h33b == _GEN_7426 ? ram_827 : _GEN_826; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_828 = 10'h33c == _GEN_7426 ? ram_828 : _GEN_827; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_829 = 10'h33d == _GEN_7426 ? ram_829 : _GEN_828; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_830 = 10'h33e == _GEN_7426 ? ram_830 : _GEN_829; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_831 = 10'h33f == _GEN_7426 ? ram_831 : _GEN_830; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_832 = 10'h340 == _GEN_7426 ? ram_832 : _GEN_831; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_833 = 10'h341 == _GEN_7426 ? ram_833 : _GEN_832; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_834 = 10'h342 == _GEN_7426 ? ram_834 : _GEN_833; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_835 = 10'h343 == _GEN_7426 ? ram_835 : _GEN_834; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_836 = 10'h344 == _GEN_7426 ? ram_836 : _GEN_835; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_837 = 10'h345 == _GEN_7426 ? ram_837 : _GEN_836; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_838 = 10'h346 == _GEN_7426 ? ram_838 : _GEN_837; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_839 = 10'h347 == _GEN_7426 ? ram_839 : _GEN_838; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_840 = 10'h348 == _GEN_7426 ? ram_840 : _GEN_839; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_841 = 10'h349 == _GEN_7426 ? ram_841 : _GEN_840; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_842 = 10'h34a == _GEN_7426 ? ram_842 : _GEN_841; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_843 = 10'h34b == _GEN_7426 ? ram_843 : _GEN_842; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_844 = 10'h34c == _GEN_7426 ? ram_844 : _GEN_843; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_845 = 10'h34d == _GEN_7426 ? ram_845 : _GEN_844; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_846 = 10'h34e == _GEN_7426 ? ram_846 : _GEN_845; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_847 = 10'h34f == _GEN_7426 ? ram_847 : _GEN_846; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_848 = 10'h350 == _GEN_7426 ? ram_848 : _GEN_847; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_849 = 10'h351 == _GEN_7426 ? ram_849 : _GEN_848; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_850 = 10'h352 == _GEN_7426 ? ram_850 : _GEN_849; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_851 = 10'h353 == _GEN_7426 ? ram_851 : _GEN_850; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_852 = 10'h354 == _GEN_7426 ? ram_852 : _GEN_851; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_853 = 10'h355 == _GEN_7426 ? ram_853 : _GEN_852; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_854 = 10'h356 == _GEN_7426 ? ram_854 : _GEN_853; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_855 = 10'h357 == _GEN_7426 ? ram_855 : _GEN_854; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_856 = 10'h358 == _GEN_7426 ? ram_856 : _GEN_855; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_857 = 10'h359 == _GEN_7426 ? ram_857 : _GEN_856; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_858 = 10'h35a == _GEN_7426 ? ram_858 : _GEN_857; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_859 = 10'h35b == _GEN_7426 ? ram_859 : _GEN_858; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_860 = 10'h35c == _GEN_7426 ? ram_860 : _GEN_859; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_861 = 10'h35d == _GEN_7426 ? ram_861 : _GEN_860; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_862 = 10'h35e == _GEN_7426 ? ram_862 : _GEN_861; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_863 = 10'h35f == _GEN_7426 ? ram_863 : _GEN_862; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_864 = 10'h360 == _GEN_7426 ? ram_864 : _GEN_863; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_865 = 10'h361 == _GEN_7426 ? ram_865 : _GEN_864; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_866 = 10'h362 == _GEN_7426 ? ram_866 : _GEN_865; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_867 = 10'h363 == _GEN_7426 ? ram_867 : _GEN_866; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_868 = 10'h364 == _GEN_7426 ? ram_868 : _GEN_867; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_869 = 10'h365 == _GEN_7426 ? ram_869 : _GEN_868; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_870 = 10'h366 == _GEN_7426 ? ram_870 : _GEN_869; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_871 = 10'h367 == _GEN_7426 ? ram_871 : _GEN_870; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_872 = 10'h368 == _GEN_7426 ? ram_872 : _GEN_871; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_873 = 10'h369 == _GEN_7426 ? ram_873 : _GEN_872; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_874 = 10'h36a == _GEN_7426 ? ram_874 : _GEN_873; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_875 = 10'h36b == _GEN_7426 ? ram_875 : _GEN_874; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_876 = 10'h36c == _GEN_7426 ? ram_876 : _GEN_875; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_877 = 10'h36d == _GEN_7426 ? ram_877 : _GEN_876; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_878 = 10'h36e == _GEN_7426 ? ram_878 : _GEN_877; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_879 = 10'h36f == _GEN_7426 ? ram_879 : _GEN_878; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_880 = 10'h370 == _GEN_7426 ? ram_880 : _GEN_879; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_881 = 10'h371 == _GEN_7426 ? ram_881 : _GEN_880; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_882 = 10'h372 == _GEN_7426 ? ram_882 : _GEN_881; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_883 = 10'h373 == _GEN_7426 ? ram_883 : _GEN_882; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_884 = 10'h374 == _GEN_7426 ? ram_884 : _GEN_883; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_885 = 10'h375 == _GEN_7426 ? ram_885 : _GEN_884; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_886 = 10'h376 == _GEN_7426 ? ram_886 : _GEN_885; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_887 = 10'h377 == _GEN_7426 ? ram_887 : _GEN_886; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_888 = 10'h378 == _GEN_7426 ? ram_888 : _GEN_887; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_889 = 10'h379 == _GEN_7426 ? ram_889 : _GEN_888; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_890 = 10'h37a == _GEN_7426 ? ram_890 : _GEN_889; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_891 = 10'h37b == _GEN_7426 ? ram_891 : _GEN_890; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_892 = 10'h37c == _GEN_7426 ? ram_892 : _GEN_891; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_893 = 10'h37d == _GEN_7426 ? ram_893 : _GEN_892; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_894 = 10'h37e == _GEN_7426 ? ram_894 : _GEN_893; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_895 = 10'h37f == _GEN_7426 ? ram_895 : _GEN_894; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_896 = 10'h380 == _GEN_7426 ? ram_896 : _GEN_895; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_897 = 10'h381 == _GEN_7426 ? ram_897 : _GEN_896; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_898 = 10'h382 == _GEN_7426 ? ram_898 : _GEN_897; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_899 = 10'h383 == _GEN_7426 ? ram_899 : _GEN_898; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_900 = 10'h384 == _GEN_7426 ? ram_900 : _GEN_899; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_901 = 10'h385 == _GEN_7426 ? ram_901 : _GEN_900; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_902 = 10'h386 == _GEN_7426 ? ram_902 : _GEN_901; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_903 = 10'h387 == _GEN_7426 ? ram_903 : _GEN_902; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_904 = 10'h388 == _GEN_7426 ? ram_904 : _GEN_903; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_905 = 10'h389 == _GEN_7426 ? ram_905 : _GEN_904; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_906 = 10'h38a == _GEN_7426 ? ram_906 : _GEN_905; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_907 = 10'h38b == _GEN_7426 ? ram_907 : _GEN_906; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_908 = 10'h38c == _GEN_7426 ? ram_908 : _GEN_907; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_909 = 10'h38d == _GEN_7426 ? ram_909 : _GEN_908; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_910 = 10'h38e == _GEN_7426 ? ram_910 : _GEN_909; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_911 = 10'h38f == _GEN_7426 ? ram_911 : _GEN_910; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_912 = 10'h390 == _GEN_7426 ? ram_912 : _GEN_911; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_913 = 10'h391 == _GEN_7426 ? ram_913 : _GEN_912; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_914 = 10'h392 == _GEN_7426 ? ram_914 : _GEN_913; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_915 = 10'h393 == _GEN_7426 ? ram_915 : _GEN_914; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_916 = 10'h394 == _GEN_7426 ? ram_916 : _GEN_915; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_917 = 10'h395 == _GEN_7426 ? ram_917 : _GEN_916; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_918 = 10'h396 == _GEN_7426 ? ram_918 : _GEN_917; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_919 = 10'h397 == _GEN_7426 ? ram_919 : _GEN_918; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_920 = 10'h398 == _GEN_7426 ? ram_920 : _GEN_919; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_921 = 10'h399 == _GEN_7426 ? ram_921 : _GEN_920; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_922 = 10'h39a == _GEN_7426 ? ram_922 : _GEN_921; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_923 = 10'h39b == _GEN_7426 ? ram_923 : _GEN_922; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_924 = 10'h39c == _GEN_7426 ? ram_924 : _GEN_923; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_925 = 10'h39d == _GEN_7426 ? ram_925 : _GEN_924; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_926 = 10'h39e == _GEN_7426 ? ram_926 : _GEN_925; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_927 = 10'h39f == _GEN_7426 ? ram_927 : _GEN_926; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_928 = 10'h3a0 == _GEN_7426 ? ram_928 : _GEN_927; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_929 = 10'h3a1 == _GEN_7426 ? ram_929 : _GEN_928; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_930 = 10'h3a2 == _GEN_7426 ? ram_930 : _GEN_929; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_931 = 10'h3a3 == _GEN_7426 ? ram_931 : _GEN_930; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_932 = 10'h3a4 == _GEN_7426 ? ram_932 : _GEN_931; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_933 = 10'h3a5 == _GEN_7426 ? ram_933 : _GEN_932; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_934 = 10'h3a6 == _GEN_7426 ? ram_934 : _GEN_933; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_935 = 10'h3a7 == _GEN_7426 ? ram_935 : _GEN_934; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_936 = 10'h3a8 == _GEN_7426 ? ram_936 : _GEN_935; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_937 = 10'h3a9 == _GEN_7426 ? ram_937 : _GEN_936; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_938 = 10'h3aa == _GEN_7426 ? ram_938 : _GEN_937; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_939 = 10'h3ab == _GEN_7426 ? ram_939 : _GEN_938; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_940 = 10'h3ac == _GEN_7426 ? ram_940 : _GEN_939; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_941 = 10'h3ad == _GEN_7426 ? ram_941 : _GEN_940; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_942 = 10'h3ae == _GEN_7426 ? ram_942 : _GEN_941; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_943 = 10'h3af == _GEN_7426 ? ram_943 : _GEN_942; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_944 = 10'h3b0 == _GEN_7426 ? ram_944 : _GEN_943; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_945 = 10'h3b1 == _GEN_7426 ? ram_945 : _GEN_944; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_946 = 10'h3b2 == _GEN_7426 ? ram_946 : _GEN_945; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_947 = 10'h3b3 == _GEN_7426 ? ram_947 : _GEN_946; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_948 = 10'h3b4 == _GEN_7426 ? ram_948 : _GEN_947; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_949 = 10'h3b5 == _GEN_7426 ? ram_949 : _GEN_948; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_950 = 10'h3b6 == _GEN_7426 ? ram_950 : _GEN_949; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_951 = 10'h3b7 == _GEN_7426 ? ram_951 : _GEN_950; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_952 = 10'h3b8 == _GEN_7426 ? ram_952 : _GEN_951; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_953 = 10'h3b9 == _GEN_7426 ? ram_953 : _GEN_952; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_954 = 10'h3ba == _GEN_7426 ? ram_954 : _GEN_953; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_955 = 10'h3bb == _GEN_7426 ? ram_955 : _GEN_954; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_956 = 10'h3bc == _GEN_7426 ? ram_956 : _GEN_955; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_957 = 10'h3bd == _GEN_7426 ? ram_957 : _GEN_956; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_958 = 10'h3be == _GEN_7426 ? ram_958 : _GEN_957; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_959 = 10'h3bf == _GEN_7426 ? ram_959 : _GEN_958; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_960 = 10'h3c0 == _GEN_7426 ? ram_960 : _GEN_959; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_961 = 10'h3c1 == _GEN_7426 ? ram_961 : _GEN_960; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_962 = 10'h3c2 == _GEN_7426 ? ram_962 : _GEN_961; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_963 = 10'h3c3 == _GEN_7426 ? ram_963 : _GEN_962; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_964 = 10'h3c4 == _GEN_7426 ? ram_964 : _GEN_963; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_965 = 10'h3c5 == _GEN_7426 ? ram_965 : _GEN_964; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_966 = 10'h3c6 == _GEN_7426 ? ram_966 : _GEN_965; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_967 = 10'h3c7 == _GEN_7426 ? ram_967 : _GEN_966; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_968 = 10'h3c8 == _GEN_7426 ? ram_968 : _GEN_967; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_969 = 10'h3c9 == _GEN_7426 ? ram_969 : _GEN_968; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_970 = 10'h3ca == _GEN_7426 ? ram_970 : _GEN_969; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_971 = 10'h3cb == _GEN_7426 ? ram_971 : _GEN_970; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_972 = 10'h3cc == _GEN_7426 ? ram_972 : _GEN_971; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_973 = 10'h3cd == _GEN_7426 ? ram_973 : _GEN_972; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_974 = 10'h3ce == _GEN_7426 ? ram_974 : _GEN_973; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_975 = 10'h3cf == _GEN_7426 ? ram_975 : _GEN_974; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_976 = 10'h3d0 == _GEN_7426 ? ram_976 : _GEN_975; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_977 = 10'h3d1 == _GEN_7426 ? ram_977 : _GEN_976; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_978 = 10'h3d2 == _GEN_7426 ? ram_978 : _GEN_977; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_979 = 10'h3d3 == _GEN_7426 ? ram_979 : _GEN_978; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_980 = 10'h3d4 == _GEN_7426 ? ram_980 : _GEN_979; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_981 = 10'h3d5 == _GEN_7426 ? ram_981 : _GEN_980; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_982 = 10'h3d6 == _GEN_7426 ? ram_982 : _GEN_981; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_983 = 10'h3d7 == _GEN_7426 ? ram_983 : _GEN_982; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_984 = 10'h3d8 == _GEN_7426 ? ram_984 : _GEN_983; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_985 = 10'h3d9 == _GEN_7426 ? ram_985 : _GEN_984; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_986 = 10'h3da == _GEN_7426 ? ram_986 : _GEN_985; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_987 = 10'h3db == _GEN_7426 ? ram_987 : _GEN_986; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_988 = 10'h3dc == _GEN_7426 ? ram_988 : _GEN_987; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_989 = 10'h3dd == _GEN_7426 ? ram_989 : _GEN_988; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_990 = 10'h3de == _GEN_7426 ? ram_990 : _GEN_989; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_991 = 10'h3df == _GEN_7426 ? ram_991 : _GEN_990; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_992 = 10'h3e0 == _GEN_7426 ? ram_992 : _GEN_991; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_993 = 10'h3e1 == _GEN_7426 ? ram_993 : _GEN_992; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_994 = 10'h3e2 == _GEN_7426 ? ram_994 : _GEN_993; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_995 = 10'h3e3 == _GEN_7426 ? ram_995 : _GEN_994; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_996 = 10'h3e4 == _GEN_7426 ? ram_996 : _GEN_995; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_997 = 10'h3e5 == _GEN_7426 ? ram_997 : _GEN_996; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_998 = 10'h3e6 == _GEN_7426 ? ram_998 : _GEN_997; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_999 = 10'h3e7 == _GEN_7426 ? ram_999 : _GEN_998; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1000 = 10'h3e8 == _GEN_7426 ? ram_1000 : _GEN_999; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1001 = 10'h3e9 == _GEN_7426 ? ram_1001 : _GEN_1000; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1002 = 10'h3ea == _GEN_7426 ? ram_1002 : _GEN_1001; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1003 = 10'h3eb == _GEN_7426 ? ram_1003 : _GEN_1002; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1004 = 10'h3ec == _GEN_7426 ? ram_1004 : _GEN_1003; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1005 = 10'h3ed == _GEN_7426 ? ram_1005 : _GEN_1004; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1006 = 10'h3ee == _GEN_7426 ? ram_1006 : _GEN_1005; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1007 = 10'h3ef == _GEN_7426 ? ram_1007 : _GEN_1006; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1008 = 10'h3f0 == _GEN_7426 ? ram_1008 : _GEN_1007; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1009 = 10'h3f1 == _GEN_7426 ? ram_1009 : _GEN_1008; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1010 = 10'h3f2 == _GEN_7426 ? ram_1010 : _GEN_1009; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1011 = 10'h3f3 == _GEN_7426 ? ram_1011 : _GEN_1010; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1012 = 10'h3f4 == _GEN_7426 ? ram_1012 : _GEN_1011; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1013 = 10'h3f5 == _GEN_7426 ? ram_1013 : _GEN_1012; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1014 = 10'h3f6 == _GEN_7426 ? ram_1014 : _GEN_1013; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1015 = 10'h3f7 == _GEN_7426 ? ram_1015 : _GEN_1014; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1016 = 10'h3f8 == _GEN_7426 ? ram_1016 : _GEN_1015; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1017 = 10'h3f9 == _GEN_7426 ? ram_1017 : _GEN_1016; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1018 = 10'h3fa == _GEN_7426 ? ram_1018 : _GEN_1017; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1019 = 10'h3fb == _GEN_7426 ? ram_1019 : _GEN_1018; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1020 = 10'h3fc == _GEN_7426 ? ram_1020 : _GEN_1019; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1021 = 10'h3fd == _GEN_7426 ? ram_1021 : _GEN_1020; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1022 = 10'h3fe == _GEN_7426 ? ram_1022 : _GEN_1021; // @[DataMemory.scala 42:{28,28}]
  wire [31:0] _GEN_1023 = 10'h3ff == _GEN_7426 ? ram_1023 : _GEN_1022; // @[DataMemory.scala 42:{28,28}]
  wire [7:0] _io_readData_T_6 = 2'h1 == io_addr[1:0] ? _GEN_1023[15:8] : _GEN_1023[7:0]; // @[Mux.scala 81:58]
  wire [7:0] _io_readData_T_8 = 2'h2 == io_addr[1:0] ? _GEN_1023[23:16] : _io_readData_T_6; // @[Mux.scala 81:58]
  wire [7:0] _io_readData_T_10 = 2'h3 == io_addr[1:0] ? _GEN_1023[31:24] : _io_readData_T_8; // @[Mux.scala 81:58]
  wire [8:0] _io_readData_T_11 = {1'h0,_io_readData_T_10}; // @[Cat.scala 31:58]
  wire [7:0] bData = io_writeData[7:0]; // @[DataMemory.scala 66:31]
  wire [31:0] _ram_T_2 = {_GEN_1023[31:8],bData}; // @[Cat.scala 31:58]
  wire [31:0] _ram_T_5 = {_GEN_1023[31:16],bData,_GEN_1023[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _ram_T_8 = {_GEN_1023[31:24],bData,_GEN_1023[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _ram_T_10 = {bData,_GEN_1023[23:0]}; // @[Cat.scala 31:58]
  wire [31:0] _ram_T_12 = 2'h1 == io_addr[1:0] ? _ram_T_5 : _ram_T_2; // @[Mux.scala 81:58]
  wire [31:0] _ram_T_14 = 2'h2 == io_addr[1:0] ? _ram_T_8 : _ram_T_12; // @[Mux.scala 81:58]
  assign io_readData = {{23'd0}, _io_readData_T_11}; // @[DataMemory.scala 34:29 35:17]
  always @(posedge clock) begin
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_0 <= 32'h6c6c6548; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h0 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_0 <= _ram_T_10;
        end else begin
          ram_0 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1 <= 32'h77202c6f; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h1 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1 <= _ram_T_10;
        end else begin
          ram_1 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_2 <= 32'h646c726f; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h2 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_2 <= _ram_T_10;
        end else begin
          ram_2 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_3 <= 32'ha21; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h3 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_3 <= _ram_T_10;
        end else begin
          ram_3 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_4 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h4 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_4 <= _ram_T_10;
        end else begin
          ram_4 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_5 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h5 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_5 <= _ram_T_10;
        end else begin
          ram_5 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_6 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h6 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_6 <= _ram_T_10;
        end else begin
          ram_6 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_7 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h7 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_7 <= _ram_T_10;
        end else begin
          ram_7 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_8 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h8 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_8 <= _ram_T_10;
        end else begin
          ram_8 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_9 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h9 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_9 <= _ram_T_10;
        end else begin
          ram_9 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_10 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_10 <= _ram_T_10;
        end else begin
          ram_10 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_11 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_11 <= _ram_T_10;
        end else begin
          ram_11 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_12 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_12 <= _ram_T_10;
        end else begin
          ram_12 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_13 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_13 <= _ram_T_10;
        end else begin
          ram_13 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_14 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_14 <= _ram_T_10;
        end else begin
          ram_14 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_15 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_15 <= _ram_T_10;
        end else begin
          ram_15 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_16 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h10 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_16 <= _ram_T_10;
        end else begin
          ram_16 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_17 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h11 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_17 <= _ram_T_10;
        end else begin
          ram_17 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_18 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h12 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_18 <= _ram_T_10;
        end else begin
          ram_18 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_19 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h13 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_19 <= _ram_T_10;
        end else begin
          ram_19 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_20 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h14 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_20 <= _ram_T_10;
        end else begin
          ram_20 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_21 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h15 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_21 <= _ram_T_10;
        end else begin
          ram_21 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_22 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h16 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_22 <= _ram_T_10;
        end else begin
          ram_22 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_23 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h17 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_23 <= _ram_T_10;
        end else begin
          ram_23 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_24 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h18 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_24 <= _ram_T_10;
        end else begin
          ram_24 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_25 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h19 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_25 <= _ram_T_10;
        end else begin
          ram_25 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_26 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h1a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_26 <= _ram_T_10;
        end else begin
          ram_26 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_27 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h1b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_27 <= _ram_T_10;
        end else begin
          ram_27 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_28 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h1c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_28 <= _ram_T_10;
        end else begin
          ram_28 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_29 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h1d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_29 <= _ram_T_10;
        end else begin
          ram_29 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_30 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h1e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_30 <= _ram_T_10;
        end else begin
          ram_30 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_31 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h1f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_31 <= _ram_T_10;
        end else begin
          ram_31 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_32 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h20 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_32 <= _ram_T_10;
        end else begin
          ram_32 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_33 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h21 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_33 <= _ram_T_10;
        end else begin
          ram_33 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_34 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h22 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_34 <= _ram_T_10;
        end else begin
          ram_34 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_35 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h23 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_35 <= _ram_T_10;
        end else begin
          ram_35 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_36 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h24 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_36 <= _ram_T_10;
        end else begin
          ram_36 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_37 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h25 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_37 <= _ram_T_10;
        end else begin
          ram_37 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_38 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h26 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_38 <= _ram_T_10;
        end else begin
          ram_38 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_39 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h27 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_39 <= _ram_T_10;
        end else begin
          ram_39 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_40 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h28 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_40 <= _ram_T_10;
        end else begin
          ram_40 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_41 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h29 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_41 <= _ram_T_10;
        end else begin
          ram_41 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_42 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h2a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_42 <= _ram_T_10;
        end else begin
          ram_42 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_43 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h2b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_43 <= _ram_T_10;
        end else begin
          ram_43 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_44 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h2c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_44 <= _ram_T_10;
        end else begin
          ram_44 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_45 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h2d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_45 <= _ram_T_10;
        end else begin
          ram_45 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_46 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h2e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_46 <= _ram_T_10;
        end else begin
          ram_46 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_47 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h2f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_47 <= _ram_T_10;
        end else begin
          ram_47 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_48 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h30 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_48 <= _ram_T_10;
        end else begin
          ram_48 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_49 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h31 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_49 <= _ram_T_10;
        end else begin
          ram_49 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_50 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h32 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_50 <= _ram_T_10;
        end else begin
          ram_50 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_51 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h33 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_51 <= _ram_T_10;
        end else begin
          ram_51 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_52 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h34 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_52 <= _ram_T_10;
        end else begin
          ram_52 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_53 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h35 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_53 <= _ram_T_10;
        end else begin
          ram_53 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_54 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h36 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_54 <= _ram_T_10;
        end else begin
          ram_54 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_55 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h37 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_55 <= _ram_T_10;
        end else begin
          ram_55 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_56 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h38 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_56 <= _ram_T_10;
        end else begin
          ram_56 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_57 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h39 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_57 <= _ram_T_10;
        end else begin
          ram_57 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_58 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h3a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_58 <= _ram_T_10;
        end else begin
          ram_58 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_59 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h3b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_59 <= _ram_T_10;
        end else begin
          ram_59 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_60 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h3c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_60 <= _ram_T_10;
        end else begin
          ram_60 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_61 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h3d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_61 <= _ram_T_10;
        end else begin
          ram_61 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_62 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h3e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_62 <= _ram_T_10;
        end else begin
          ram_62 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_63 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h3f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_63 <= _ram_T_10;
        end else begin
          ram_63 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_64 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h40 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_64 <= _ram_T_10;
        end else begin
          ram_64 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_65 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h41 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_65 <= _ram_T_10;
        end else begin
          ram_65 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_66 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h42 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_66 <= _ram_T_10;
        end else begin
          ram_66 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_67 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h43 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_67 <= _ram_T_10;
        end else begin
          ram_67 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_68 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h44 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_68 <= _ram_T_10;
        end else begin
          ram_68 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_69 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h45 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_69 <= _ram_T_10;
        end else begin
          ram_69 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_70 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h46 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_70 <= _ram_T_10;
        end else begin
          ram_70 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_71 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h47 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_71 <= _ram_T_10;
        end else begin
          ram_71 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_72 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h48 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_72 <= _ram_T_10;
        end else begin
          ram_72 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_73 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h49 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_73 <= _ram_T_10;
        end else begin
          ram_73 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_74 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h4a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_74 <= _ram_T_10;
        end else begin
          ram_74 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_75 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h4b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_75 <= _ram_T_10;
        end else begin
          ram_75 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_76 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h4c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_76 <= _ram_T_10;
        end else begin
          ram_76 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_77 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h4d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_77 <= _ram_T_10;
        end else begin
          ram_77 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_78 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h4e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_78 <= _ram_T_10;
        end else begin
          ram_78 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_79 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h4f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_79 <= _ram_T_10;
        end else begin
          ram_79 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_80 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h50 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_80 <= _ram_T_10;
        end else begin
          ram_80 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_81 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h51 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_81 <= _ram_T_10;
        end else begin
          ram_81 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_82 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h52 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_82 <= _ram_T_10;
        end else begin
          ram_82 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_83 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h53 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_83 <= _ram_T_10;
        end else begin
          ram_83 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_84 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h54 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_84 <= _ram_T_10;
        end else begin
          ram_84 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_85 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h55 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_85 <= _ram_T_10;
        end else begin
          ram_85 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_86 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h56 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_86 <= _ram_T_10;
        end else begin
          ram_86 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_87 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h57 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_87 <= _ram_T_10;
        end else begin
          ram_87 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_88 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h58 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_88 <= _ram_T_10;
        end else begin
          ram_88 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_89 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h59 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_89 <= _ram_T_10;
        end else begin
          ram_89 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_90 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h5a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_90 <= _ram_T_10;
        end else begin
          ram_90 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_91 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h5b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_91 <= _ram_T_10;
        end else begin
          ram_91 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_92 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h5c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_92 <= _ram_T_10;
        end else begin
          ram_92 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_93 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h5d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_93 <= _ram_T_10;
        end else begin
          ram_93 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_94 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h5e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_94 <= _ram_T_10;
        end else begin
          ram_94 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_95 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h5f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_95 <= _ram_T_10;
        end else begin
          ram_95 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_96 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h60 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_96 <= _ram_T_10;
        end else begin
          ram_96 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_97 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h61 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_97 <= _ram_T_10;
        end else begin
          ram_97 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_98 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h62 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_98 <= _ram_T_10;
        end else begin
          ram_98 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_99 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h63 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_99 <= _ram_T_10;
        end else begin
          ram_99 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_100 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h64 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_100 <= _ram_T_10;
        end else begin
          ram_100 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_101 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h65 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_101 <= _ram_T_10;
        end else begin
          ram_101 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_102 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h66 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_102 <= _ram_T_10;
        end else begin
          ram_102 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_103 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h67 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_103 <= _ram_T_10;
        end else begin
          ram_103 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_104 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h68 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_104 <= _ram_T_10;
        end else begin
          ram_104 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_105 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h69 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_105 <= _ram_T_10;
        end else begin
          ram_105 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_106 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h6a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_106 <= _ram_T_10;
        end else begin
          ram_106 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_107 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h6b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_107 <= _ram_T_10;
        end else begin
          ram_107 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_108 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h6c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_108 <= _ram_T_10;
        end else begin
          ram_108 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_109 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h6d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_109 <= _ram_T_10;
        end else begin
          ram_109 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_110 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h6e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_110 <= _ram_T_10;
        end else begin
          ram_110 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_111 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h6f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_111 <= _ram_T_10;
        end else begin
          ram_111 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_112 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h70 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_112 <= _ram_T_10;
        end else begin
          ram_112 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_113 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h71 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_113 <= _ram_T_10;
        end else begin
          ram_113 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_114 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h72 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_114 <= _ram_T_10;
        end else begin
          ram_114 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_115 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h73 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_115 <= _ram_T_10;
        end else begin
          ram_115 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_116 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h74 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_116 <= _ram_T_10;
        end else begin
          ram_116 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_117 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h75 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_117 <= _ram_T_10;
        end else begin
          ram_117 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_118 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h76 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_118 <= _ram_T_10;
        end else begin
          ram_118 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_119 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h77 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_119 <= _ram_T_10;
        end else begin
          ram_119 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_120 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h78 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_120 <= _ram_T_10;
        end else begin
          ram_120 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_121 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h79 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_121 <= _ram_T_10;
        end else begin
          ram_121 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_122 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h7a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_122 <= _ram_T_10;
        end else begin
          ram_122 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_123 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h7b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_123 <= _ram_T_10;
        end else begin
          ram_123 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_124 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h7c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_124 <= _ram_T_10;
        end else begin
          ram_124 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_125 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h7d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_125 <= _ram_T_10;
        end else begin
          ram_125 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_126 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h7e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_126 <= _ram_T_10;
        end else begin
          ram_126 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_127 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h7f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_127 <= _ram_T_10;
        end else begin
          ram_127 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_128 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h80 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_128 <= _ram_T_10;
        end else begin
          ram_128 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_129 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h81 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_129 <= _ram_T_10;
        end else begin
          ram_129 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_130 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h82 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_130 <= _ram_T_10;
        end else begin
          ram_130 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_131 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h83 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_131 <= _ram_T_10;
        end else begin
          ram_131 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_132 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h84 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_132 <= _ram_T_10;
        end else begin
          ram_132 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_133 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h85 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_133 <= _ram_T_10;
        end else begin
          ram_133 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_134 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h86 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_134 <= _ram_T_10;
        end else begin
          ram_134 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_135 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h87 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_135 <= _ram_T_10;
        end else begin
          ram_135 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_136 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h88 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_136 <= _ram_T_10;
        end else begin
          ram_136 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_137 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h89 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_137 <= _ram_T_10;
        end else begin
          ram_137 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_138 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h8a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_138 <= _ram_T_10;
        end else begin
          ram_138 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_139 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h8b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_139 <= _ram_T_10;
        end else begin
          ram_139 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_140 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h8c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_140 <= _ram_T_10;
        end else begin
          ram_140 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_141 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h8d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_141 <= _ram_T_10;
        end else begin
          ram_141 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_142 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h8e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_142 <= _ram_T_10;
        end else begin
          ram_142 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_143 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h8f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_143 <= _ram_T_10;
        end else begin
          ram_143 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_144 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h90 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_144 <= _ram_T_10;
        end else begin
          ram_144 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_145 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h91 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_145 <= _ram_T_10;
        end else begin
          ram_145 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_146 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h92 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_146 <= _ram_T_10;
        end else begin
          ram_146 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_147 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h93 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_147 <= _ram_T_10;
        end else begin
          ram_147 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_148 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h94 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_148 <= _ram_T_10;
        end else begin
          ram_148 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_149 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h95 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_149 <= _ram_T_10;
        end else begin
          ram_149 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_150 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h96 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_150 <= _ram_T_10;
        end else begin
          ram_150 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_151 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h97 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_151 <= _ram_T_10;
        end else begin
          ram_151 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_152 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h98 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_152 <= _ram_T_10;
        end else begin
          ram_152 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_153 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h99 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_153 <= _ram_T_10;
        end else begin
          ram_153 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_154 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h9a == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_154 <= _ram_T_10;
        end else begin
          ram_154 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_155 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h9b == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_155 <= _ram_T_10;
        end else begin
          ram_155 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_156 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h9c == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_156 <= _ram_T_10;
        end else begin
          ram_156 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_157 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h9d == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_157 <= _ram_T_10;
        end else begin
          ram_157 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_158 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h9e == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_158 <= _ram_T_10;
        end else begin
          ram_158 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_159 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'h9f == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_159 <= _ram_T_10;
        end else begin
          ram_159 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_160 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha0 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_160 <= _ram_T_10;
        end else begin
          ram_160 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_161 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha1 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_161 <= _ram_T_10;
        end else begin
          ram_161 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_162 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha2 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_162 <= _ram_T_10;
        end else begin
          ram_162 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_163 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha3 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_163 <= _ram_T_10;
        end else begin
          ram_163 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_164 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha4 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_164 <= _ram_T_10;
        end else begin
          ram_164 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_165 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha5 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_165 <= _ram_T_10;
        end else begin
          ram_165 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_166 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha6 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_166 <= _ram_T_10;
        end else begin
          ram_166 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_167 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha7 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_167 <= _ram_T_10;
        end else begin
          ram_167 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_168 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha8 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_168 <= _ram_T_10;
        end else begin
          ram_168 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_169 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'ha9 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_169 <= _ram_T_10;
        end else begin
          ram_169 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_170 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'haa == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_170 <= _ram_T_10;
        end else begin
          ram_170 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_171 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hab == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_171 <= _ram_T_10;
        end else begin
          ram_171 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_172 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hac == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_172 <= _ram_T_10;
        end else begin
          ram_172 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_173 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'had == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_173 <= _ram_T_10;
        end else begin
          ram_173 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_174 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hae == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_174 <= _ram_T_10;
        end else begin
          ram_174 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_175 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'haf == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_175 <= _ram_T_10;
        end else begin
          ram_175 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_176 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb0 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_176 <= _ram_T_10;
        end else begin
          ram_176 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_177 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb1 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_177 <= _ram_T_10;
        end else begin
          ram_177 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_178 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb2 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_178 <= _ram_T_10;
        end else begin
          ram_178 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_179 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb3 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_179 <= _ram_T_10;
        end else begin
          ram_179 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_180 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb4 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_180 <= _ram_T_10;
        end else begin
          ram_180 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_181 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb5 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_181 <= _ram_T_10;
        end else begin
          ram_181 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_182 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb6 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_182 <= _ram_T_10;
        end else begin
          ram_182 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_183 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb7 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_183 <= _ram_T_10;
        end else begin
          ram_183 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_184 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb8 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_184 <= _ram_T_10;
        end else begin
          ram_184 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_185 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hb9 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_185 <= _ram_T_10;
        end else begin
          ram_185 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_186 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hba == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_186 <= _ram_T_10;
        end else begin
          ram_186 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_187 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hbb == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_187 <= _ram_T_10;
        end else begin
          ram_187 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_188 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hbc == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_188 <= _ram_T_10;
        end else begin
          ram_188 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_189 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hbd == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_189 <= _ram_T_10;
        end else begin
          ram_189 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_190 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hbe == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_190 <= _ram_T_10;
        end else begin
          ram_190 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_191 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hbf == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_191 <= _ram_T_10;
        end else begin
          ram_191 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_192 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc0 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_192 <= _ram_T_10;
        end else begin
          ram_192 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_193 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc1 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_193 <= _ram_T_10;
        end else begin
          ram_193 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_194 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc2 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_194 <= _ram_T_10;
        end else begin
          ram_194 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_195 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc3 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_195 <= _ram_T_10;
        end else begin
          ram_195 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_196 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc4 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_196 <= _ram_T_10;
        end else begin
          ram_196 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_197 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc5 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_197 <= _ram_T_10;
        end else begin
          ram_197 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_198 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc6 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_198 <= _ram_T_10;
        end else begin
          ram_198 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_199 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc7 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_199 <= _ram_T_10;
        end else begin
          ram_199 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_200 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc8 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_200 <= _ram_T_10;
        end else begin
          ram_200 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_201 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hc9 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_201 <= _ram_T_10;
        end else begin
          ram_201 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_202 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hca == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_202 <= _ram_T_10;
        end else begin
          ram_202 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_203 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hcb == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_203 <= _ram_T_10;
        end else begin
          ram_203 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_204 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hcc == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_204 <= _ram_T_10;
        end else begin
          ram_204 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_205 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hcd == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_205 <= _ram_T_10;
        end else begin
          ram_205 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_206 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hce == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_206 <= _ram_T_10;
        end else begin
          ram_206 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_207 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hcf == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_207 <= _ram_T_10;
        end else begin
          ram_207 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_208 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd0 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_208 <= _ram_T_10;
        end else begin
          ram_208 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_209 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd1 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_209 <= _ram_T_10;
        end else begin
          ram_209 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_210 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd2 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_210 <= _ram_T_10;
        end else begin
          ram_210 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_211 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd3 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_211 <= _ram_T_10;
        end else begin
          ram_211 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_212 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd4 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_212 <= _ram_T_10;
        end else begin
          ram_212 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_213 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd5 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_213 <= _ram_T_10;
        end else begin
          ram_213 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_214 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd6 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_214 <= _ram_T_10;
        end else begin
          ram_214 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_215 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd7 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_215 <= _ram_T_10;
        end else begin
          ram_215 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_216 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd8 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_216 <= _ram_T_10;
        end else begin
          ram_216 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_217 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hd9 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_217 <= _ram_T_10;
        end else begin
          ram_217 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_218 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hda == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_218 <= _ram_T_10;
        end else begin
          ram_218 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_219 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hdb == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_219 <= _ram_T_10;
        end else begin
          ram_219 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_220 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hdc == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_220 <= _ram_T_10;
        end else begin
          ram_220 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_221 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hdd == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_221 <= _ram_T_10;
        end else begin
          ram_221 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_222 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hde == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_222 <= _ram_T_10;
        end else begin
          ram_222 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_223 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hdf == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_223 <= _ram_T_10;
        end else begin
          ram_223 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_224 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he0 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_224 <= _ram_T_10;
        end else begin
          ram_224 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_225 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he1 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_225 <= _ram_T_10;
        end else begin
          ram_225 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_226 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he2 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_226 <= _ram_T_10;
        end else begin
          ram_226 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_227 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he3 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_227 <= _ram_T_10;
        end else begin
          ram_227 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_228 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he4 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_228 <= _ram_T_10;
        end else begin
          ram_228 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_229 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he5 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_229 <= _ram_T_10;
        end else begin
          ram_229 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_230 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he6 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_230 <= _ram_T_10;
        end else begin
          ram_230 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_231 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he7 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_231 <= _ram_T_10;
        end else begin
          ram_231 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_232 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he8 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_232 <= _ram_T_10;
        end else begin
          ram_232 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_233 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'he9 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_233 <= _ram_T_10;
        end else begin
          ram_233 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_234 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hea == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_234 <= _ram_T_10;
        end else begin
          ram_234 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_235 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'heb == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_235 <= _ram_T_10;
        end else begin
          ram_235 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_236 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hec == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_236 <= _ram_T_10;
        end else begin
          ram_236 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_237 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hed == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_237 <= _ram_T_10;
        end else begin
          ram_237 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_238 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hee == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_238 <= _ram_T_10;
        end else begin
          ram_238 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_239 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hef == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_239 <= _ram_T_10;
        end else begin
          ram_239 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_240 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf0 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_240 <= _ram_T_10;
        end else begin
          ram_240 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_241 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf1 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_241 <= _ram_T_10;
        end else begin
          ram_241 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_242 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf2 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_242 <= _ram_T_10;
        end else begin
          ram_242 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_243 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf3 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_243 <= _ram_T_10;
        end else begin
          ram_243 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_244 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf4 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_244 <= _ram_T_10;
        end else begin
          ram_244 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_245 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf5 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_245 <= _ram_T_10;
        end else begin
          ram_245 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_246 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf6 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_246 <= _ram_T_10;
        end else begin
          ram_246 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_247 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf7 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_247 <= _ram_T_10;
        end else begin
          ram_247 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_248 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf8 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_248 <= _ram_T_10;
        end else begin
          ram_248 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_249 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hf9 == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_249 <= _ram_T_10;
        end else begin
          ram_249 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_250 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hfa == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_250 <= _ram_T_10;
        end else begin
          ram_250 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_251 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hfb == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_251 <= _ram_T_10;
        end else begin
          ram_251 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_252 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hfc == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_252 <= _ram_T_10;
        end else begin
          ram_252 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_253 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hfd == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_253 <= _ram_T_10;
        end else begin
          ram_253 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_254 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hfe == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_254 <= _ram_T_10;
        end else begin
          ram_254 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_255 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (8'hff == io_addr[9:2]) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_255 <= _ram_T_10;
        end else begin
          ram_255 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_256 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h100 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_256 <= _ram_T_10;
        end else begin
          ram_256 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_257 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h101 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_257 <= _ram_T_10;
        end else begin
          ram_257 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_258 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h102 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_258 <= _ram_T_10;
        end else begin
          ram_258 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_259 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h103 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_259 <= _ram_T_10;
        end else begin
          ram_259 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_260 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h104 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_260 <= _ram_T_10;
        end else begin
          ram_260 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_261 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h105 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_261 <= _ram_T_10;
        end else begin
          ram_261 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_262 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h106 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_262 <= _ram_T_10;
        end else begin
          ram_262 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_263 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h107 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_263 <= _ram_T_10;
        end else begin
          ram_263 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_264 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h108 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_264 <= _ram_T_10;
        end else begin
          ram_264 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_265 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h109 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_265 <= _ram_T_10;
        end else begin
          ram_265 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_266 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h10a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_266 <= _ram_T_10;
        end else begin
          ram_266 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_267 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h10b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_267 <= _ram_T_10;
        end else begin
          ram_267 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_268 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h10c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_268 <= _ram_T_10;
        end else begin
          ram_268 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_269 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h10d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_269 <= _ram_T_10;
        end else begin
          ram_269 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_270 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h10e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_270 <= _ram_T_10;
        end else begin
          ram_270 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_271 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h10f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_271 <= _ram_T_10;
        end else begin
          ram_271 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_272 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h110 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_272 <= _ram_T_10;
        end else begin
          ram_272 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_273 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h111 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_273 <= _ram_T_10;
        end else begin
          ram_273 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_274 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h112 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_274 <= _ram_T_10;
        end else begin
          ram_274 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_275 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h113 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_275 <= _ram_T_10;
        end else begin
          ram_275 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_276 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h114 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_276 <= _ram_T_10;
        end else begin
          ram_276 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_277 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h115 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_277 <= _ram_T_10;
        end else begin
          ram_277 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_278 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h116 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_278 <= _ram_T_10;
        end else begin
          ram_278 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_279 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h117 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_279 <= _ram_T_10;
        end else begin
          ram_279 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_280 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h118 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_280 <= _ram_T_10;
        end else begin
          ram_280 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_281 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h119 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_281 <= _ram_T_10;
        end else begin
          ram_281 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_282 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h11a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_282 <= _ram_T_10;
        end else begin
          ram_282 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_283 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h11b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_283 <= _ram_T_10;
        end else begin
          ram_283 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_284 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h11c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_284 <= _ram_T_10;
        end else begin
          ram_284 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_285 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h11d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_285 <= _ram_T_10;
        end else begin
          ram_285 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_286 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h11e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_286 <= _ram_T_10;
        end else begin
          ram_286 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_287 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h11f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_287 <= _ram_T_10;
        end else begin
          ram_287 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_288 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h120 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_288 <= _ram_T_10;
        end else begin
          ram_288 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_289 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h121 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_289 <= _ram_T_10;
        end else begin
          ram_289 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_290 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h122 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_290 <= _ram_T_10;
        end else begin
          ram_290 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_291 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h123 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_291 <= _ram_T_10;
        end else begin
          ram_291 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_292 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h124 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_292 <= _ram_T_10;
        end else begin
          ram_292 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_293 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h125 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_293 <= _ram_T_10;
        end else begin
          ram_293 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_294 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h126 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_294 <= _ram_T_10;
        end else begin
          ram_294 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_295 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h127 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_295 <= _ram_T_10;
        end else begin
          ram_295 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_296 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h128 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_296 <= _ram_T_10;
        end else begin
          ram_296 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_297 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h129 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_297 <= _ram_T_10;
        end else begin
          ram_297 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_298 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h12a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_298 <= _ram_T_10;
        end else begin
          ram_298 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_299 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h12b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_299 <= _ram_T_10;
        end else begin
          ram_299 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_300 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h12c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_300 <= _ram_T_10;
        end else begin
          ram_300 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_301 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h12d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_301 <= _ram_T_10;
        end else begin
          ram_301 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_302 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h12e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_302 <= _ram_T_10;
        end else begin
          ram_302 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_303 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h12f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_303 <= _ram_T_10;
        end else begin
          ram_303 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_304 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h130 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_304 <= _ram_T_10;
        end else begin
          ram_304 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_305 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h131 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_305 <= _ram_T_10;
        end else begin
          ram_305 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_306 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h132 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_306 <= _ram_T_10;
        end else begin
          ram_306 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_307 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h133 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_307 <= _ram_T_10;
        end else begin
          ram_307 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_308 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h134 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_308 <= _ram_T_10;
        end else begin
          ram_308 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_309 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h135 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_309 <= _ram_T_10;
        end else begin
          ram_309 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_310 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h136 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_310 <= _ram_T_10;
        end else begin
          ram_310 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_311 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h137 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_311 <= _ram_T_10;
        end else begin
          ram_311 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_312 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h138 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_312 <= _ram_T_10;
        end else begin
          ram_312 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_313 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h139 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_313 <= _ram_T_10;
        end else begin
          ram_313 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_314 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h13a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_314 <= _ram_T_10;
        end else begin
          ram_314 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_315 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h13b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_315 <= _ram_T_10;
        end else begin
          ram_315 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_316 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h13c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_316 <= _ram_T_10;
        end else begin
          ram_316 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_317 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h13d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_317 <= _ram_T_10;
        end else begin
          ram_317 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_318 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h13e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_318 <= _ram_T_10;
        end else begin
          ram_318 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_319 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h13f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_319 <= _ram_T_10;
        end else begin
          ram_319 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_320 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h140 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_320 <= _ram_T_10;
        end else begin
          ram_320 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_321 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h141 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_321 <= _ram_T_10;
        end else begin
          ram_321 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_322 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h142 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_322 <= _ram_T_10;
        end else begin
          ram_322 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_323 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h143 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_323 <= _ram_T_10;
        end else begin
          ram_323 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_324 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h144 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_324 <= _ram_T_10;
        end else begin
          ram_324 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_325 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h145 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_325 <= _ram_T_10;
        end else begin
          ram_325 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_326 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h146 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_326 <= _ram_T_10;
        end else begin
          ram_326 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_327 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h147 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_327 <= _ram_T_10;
        end else begin
          ram_327 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_328 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h148 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_328 <= _ram_T_10;
        end else begin
          ram_328 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_329 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h149 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_329 <= _ram_T_10;
        end else begin
          ram_329 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_330 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h14a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_330 <= _ram_T_10;
        end else begin
          ram_330 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_331 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h14b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_331 <= _ram_T_10;
        end else begin
          ram_331 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_332 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h14c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_332 <= _ram_T_10;
        end else begin
          ram_332 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_333 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h14d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_333 <= _ram_T_10;
        end else begin
          ram_333 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_334 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h14e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_334 <= _ram_T_10;
        end else begin
          ram_334 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_335 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h14f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_335 <= _ram_T_10;
        end else begin
          ram_335 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_336 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h150 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_336 <= _ram_T_10;
        end else begin
          ram_336 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_337 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h151 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_337 <= _ram_T_10;
        end else begin
          ram_337 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_338 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h152 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_338 <= _ram_T_10;
        end else begin
          ram_338 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_339 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h153 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_339 <= _ram_T_10;
        end else begin
          ram_339 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_340 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h154 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_340 <= _ram_T_10;
        end else begin
          ram_340 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_341 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h155 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_341 <= _ram_T_10;
        end else begin
          ram_341 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_342 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h156 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_342 <= _ram_T_10;
        end else begin
          ram_342 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_343 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h157 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_343 <= _ram_T_10;
        end else begin
          ram_343 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_344 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h158 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_344 <= _ram_T_10;
        end else begin
          ram_344 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_345 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h159 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_345 <= _ram_T_10;
        end else begin
          ram_345 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_346 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h15a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_346 <= _ram_T_10;
        end else begin
          ram_346 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_347 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h15b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_347 <= _ram_T_10;
        end else begin
          ram_347 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_348 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h15c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_348 <= _ram_T_10;
        end else begin
          ram_348 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_349 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h15d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_349 <= _ram_T_10;
        end else begin
          ram_349 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_350 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h15e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_350 <= _ram_T_10;
        end else begin
          ram_350 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_351 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h15f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_351 <= _ram_T_10;
        end else begin
          ram_351 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_352 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h160 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_352 <= _ram_T_10;
        end else begin
          ram_352 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_353 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h161 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_353 <= _ram_T_10;
        end else begin
          ram_353 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_354 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h162 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_354 <= _ram_T_10;
        end else begin
          ram_354 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_355 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h163 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_355 <= _ram_T_10;
        end else begin
          ram_355 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_356 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h164 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_356 <= _ram_T_10;
        end else begin
          ram_356 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_357 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h165 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_357 <= _ram_T_10;
        end else begin
          ram_357 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_358 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h166 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_358 <= _ram_T_10;
        end else begin
          ram_358 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_359 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h167 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_359 <= _ram_T_10;
        end else begin
          ram_359 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_360 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h168 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_360 <= _ram_T_10;
        end else begin
          ram_360 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_361 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h169 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_361 <= _ram_T_10;
        end else begin
          ram_361 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_362 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h16a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_362 <= _ram_T_10;
        end else begin
          ram_362 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_363 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h16b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_363 <= _ram_T_10;
        end else begin
          ram_363 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_364 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h16c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_364 <= _ram_T_10;
        end else begin
          ram_364 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_365 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h16d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_365 <= _ram_T_10;
        end else begin
          ram_365 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_366 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h16e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_366 <= _ram_T_10;
        end else begin
          ram_366 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_367 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h16f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_367 <= _ram_T_10;
        end else begin
          ram_367 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_368 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h170 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_368 <= _ram_T_10;
        end else begin
          ram_368 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_369 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h171 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_369 <= _ram_T_10;
        end else begin
          ram_369 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_370 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h172 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_370 <= _ram_T_10;
        end else begin
          ram_370 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_371 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h173 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_371 <= _ram_T_10;
        end else begin
          ram_371 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_372 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h174 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_372 <= _ram_T_10;
        end else begin
          ram_372 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_373 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h175 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_373 <= _ram_T_10;
        end else begin
          ram_373 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_374 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h176 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_374 <= _ram_T_10;
        end else begin
          ram_374 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_375 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h177 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_375 <= _ram_T_10;
        end else begin
          ram_375 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_376 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h178 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_376 <= _ram_T_10;
        end else begin
          ram_376 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_377 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h179 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_377 <= _ram_T_10;
        end else begin
          ram_377 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_378 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h17a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_378 <= _ram_T_10;
        end else begin
          ram_378 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_379 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h17b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_379 <= _ram_T_10;
        end else begin
          ram_379 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_380 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h17c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_380 <= _ram_T_10;
        end else begin
          ram_380 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_381 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h17d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_381 <= _ram_T_10;
        end else begin
          ram_381 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_382 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h17e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_382 <= _ram_T_10;
        end else begin
          ram_382 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_383 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h17f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_383 <= _ram_T_10;
        end else begin
          ram_383 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_384 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h180 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_384 <= _ram_T_10;
        end else begin
          ram_384 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_385 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h181 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_385 <= _ram_T_10;
        end else begin
          ram_385 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_386 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h182 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_386 <= _ram_T_10;
        end else begin
          ram_386 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_387 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h183 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_387 <= _ram_T_10;
        end else begin
          ram_387 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_388 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h184 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_388 <= _ram_T_10;
        end else begin
          ram_388 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_389 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h185 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_389 <= _ram_T_10;
        end else begin
          ram_389 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_390 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h186 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_390 <= _ram_T_10;
        end else begin
          ram_390 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_391 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h187 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_391 <= _ram_T_10;
        end else begin
          ram_391 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_392 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h188 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_392 <= _ram_T_10;
        end else begin
          ram_392 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_393 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h189 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_393 <= _ram_T_10;
        end else begin
          ram_393 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_394 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h18a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_394 <= _ram_T_10;
        end else begin
          ram_394 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_395 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h18b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_395 <= _ram_T_10;
        end else begin
          ram_395 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_396 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h18c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_396 <= _ram_T_10;
        end else begin
          ram_396 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_397 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h18d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_397 <= _ram_T_10;
        end else begin
          ram_397 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_398 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h18e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_398 <= _ram_T_10;
        end else begin
          ram_398 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_399 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h18f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_399 <= _ram_T_10;
        end else begin
          ram_399 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_400 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h190 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_400 <= _ram_T_10;
        end else begin
          ram_400 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_401 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h191 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_401 <= _ram_T_10;
        end else begin
          ram_401 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_402 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h192 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_402 <= _ram_T_10;
        end else begin
          ram_402 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_403 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h193 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_403 <= _ram_T_10;
        end else begin
          ram_403 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_404 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h194 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_404 <= _ram_T_10;
        end else begin
          ram_404 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_405 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h195 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_405 <= _ram_T_10;
        end else begin
          ram_405 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_406 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h196 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_406 <= _ram_T_10;
        end else begin
          ram_406 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_407 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h197 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_407 <= _ram_T_10;
        end else begin
          ram_407 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_408 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h198 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_408 <= _ram_T_10;
        end else begin
          ram_408 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_409 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h199 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_409 <= _ram_T_10;
        end else begin
          ram_409 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_410 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h19a == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_410 <= _ram_T_10;
        end else begin
          ram_410 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_411 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h19b == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_411 <= _ram_T_10;
        end else begin
          ram_411 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_412 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h19c == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_412 <= _ram_T_10;
        end else begin
          ram_412 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_413 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h19d == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_413 <= _ram_T_10;
        end else begin
          ram_413 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_414 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h19e == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_414 <= _ram_T_10;
        end else begin
          ram_414 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_415 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h19f == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_415 <= _ram_T_10;
        end else begin
          ram_415 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_416 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a0 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_416 <= _ram_T_10;
        end else begin
          ram_416 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_417 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a1 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_417 <= _ram_T_10;
        end else begin
          ram_417 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_418 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a2 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_418 <= _ram_T_10;
        end else begin
          ram_418 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_419 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a3 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_419 <= _ram_T_10;
        end else begin
          ram_419 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_420 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a4 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_420 <= _ram_T_10;
        end else begin
          ram_420 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_421 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a5 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_421 <= _ram_T_10;
        end else begin
          ram_421 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_422 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a6 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_422 <= _ram_T_10;
        end else begin
          ram_422 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_423 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a7 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_423 <= _ram_T_10;
        end else begin
          ram_423 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_424 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a8 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_424 <= _ram_T_10;
        end else begin
          ram_424 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_425 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1a9 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_425 <= _ram_T_10;
        end else begin
          ram_425 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_426 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1aa == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_426 <= _ram_T_10;
        end else begin
          ram_426 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_427 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ab == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_427 <= _ram_T_10;
        end else begin
          ram_427 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_428 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ac == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_428 <= _ram_T_10;
        end else begin
          ram_428 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_429 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ad == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_429 <= _ram_T_10;
        end else begin
          ram_429 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_430 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ae == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_430 <= _ram_T_10;
        end else begin
          ram_430 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_431 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1af == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_431 <= _ram_T_10;
        end else begin
          ram_431 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_432 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b0 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_432 <= _ram_T_10;
        end else begin
          ram_432 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_433 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b1 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_433 <= _ram_T_10;
        end else begin
          ram_433 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_434 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b2 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_434 <= _ram_T_10;
        end else begin
          ram_434 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_435 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b3 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_435 <= _ram_T_10;
        end else begin
          ram_435 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_436 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b4 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_436 <= _ram_T_10;
        end else begin
          ram_436 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_437 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b5 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_437 <= _ram_T_10;
        end else begin
          ram_437 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_438 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b6 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_438 <= _ram_T_10;
        end else begin
          ram_438 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_439 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b7 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_439 <= _ram_T_10;
        end else begin
          ram_439 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_440 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b8 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_440 <= _ram_T_10;
        end else begin
          ram_440 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_441 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1b9 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_441 <= _ram_T_10;
        end else begin
          ram_441 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_442 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ba == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_442 <= _ram_T_10;
        end else begin
          ram_442 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_443 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1bb == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_443 <= _ram_T_10;
        end else begin
          ram_443 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_444 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1bc == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_444 <= _ram_T_10;
        end else begin
          ram_444 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_445 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1bd == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_445 <= _ram_T_10;
        end else begin
          ram_445 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_446 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1be == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_446 <= _ram_T_10;
        end else begin
          ram_446 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_447 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1bf == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_447 <= _ram_T_10;
        end else begin
          ram_447 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_448 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c0 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_448 <= _ram_T_10;
        end else begin
          ram_448 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_449 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c1 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_449 <= _ram_T_10;
        end else begin
          ram_449 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_450 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c2 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_450 <= _ram_T_10;
        end else begin
          ram_450 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_451 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c3 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_451 <= _ram_T_10;
        end else begin
          ram_451 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_452 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c4 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_452 <= _ram_T_10;
        end else begin
          ram_452 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_453 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c5 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_453 <= _ram_T_10;
        end else begin
          ram_453 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_454 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c6 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_454 <= _ram_T_10;
        end else begin
          ram_454 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_455 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c7 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_455 <= _ram_T_10;
        end else begin
          ram_455 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_456 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c8 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_456 <= _ram_T_10;
        end else begin
          ram_456 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_457 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1c9 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_457 <= _ram_T_10;
        end else begin
          ram_457 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_458 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ca == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_458 <= _ram_T_10;
        end else begin
          ram_458 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_459 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1cb == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_459 <= _ram_T_10;
        end else begin
          ram_459 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_460 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1cc == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_460 <= _ram_T_10;
        end else begin
          ram_460 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_461 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1cd == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_461 <= _ram_T_10;
        end else begin
          ram_461 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_462 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ce == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_462 <= _ram_T_10;
        end else begin
          ram_462 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_463 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1cf == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_463 <= _ram_T_10;
        end else begin
          ram_463 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_464 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d0 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_464 <= _ram_T_10;
        end else begin
          ram_464 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_465 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d1 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_465 <= _ram_T_10;
        end else begin
          ram_465 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_466 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d2 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_466 <= _ram_T_10;
        end else begin
          ram_466 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_467 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d3 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_467 <= _ram_T_10;
        end else begin
          ram_467 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_468 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d4 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_468 <= _ram_T_10;
        end else begin
          ram_468 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_469 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d5 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_469 <= _ram_T_10;
        end else begin
          ram_469 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_470 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d6 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_470 <= _ram_T_10;
        end else begin
          ram_470 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_471 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d7 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_471 <= _ram_T_10;
        end else begin
          ram_471 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_472 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d8 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_472 <= _ram_T_10;
        end else begin
          ram_472 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_473 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1d9 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_473 <= _ram_T_10;
        end else begin
          ram_473 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_474 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1da == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_474 <= _ram_T_10;
        end else begin
          ram_474 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_475 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1db == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_475 <= _ram_T_10;
        end else begin
          ram_475 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_476 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1dc == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_476 <= _ram_T_10;
        end else begin
          ram_476 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_477 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1dd == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_477 <= _ram_T_10;
        end else begin
          ram_477 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_478 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1de == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_478 <= _ram_T_10;
        end else begin
          ram_478 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_479 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1df == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_479 <= _ram_T_10;
        end else begin
          ram_479 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_480 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e0 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_480 <= _ram_T_10;
        end else begin
          ram_480 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_481 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e1 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_481 <= _ram_T_10;
        end else begin
          ram_481 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_482 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e2 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_482 <= _ram_T_10;
        end else begin
          ram_482 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_483 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e3 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_483 <= _ram_T_10;
        end else begin
          ram_483 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_484 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e4 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_484 <= _ram_T_10;
        end else begin
          ram_484 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_485 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e5 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_485 <= _ram_T_10;
        end else begin
          ram_485 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_486 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e6 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_486 <= _ram_T_10;
        end else begin
          ram_486 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_487 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e7 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_487 <= _ram_T_10;
        end else begin
          ram_487 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_488 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e8 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_488 <= _ram_T_10;
        end else begin
          ram_488 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_489 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1e9 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_489 <= _ram_T_10;
        end else begin
          ram_489 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_490 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ea == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_490 <= _ram_T_10;
        end else begin
          ram_490 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_491 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1eb == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_491 <= _ram_T_10;
        end else begin
          ram_491 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_492 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ec == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_492 <= _ram_T_10;
        end else begin
          ram_492 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_493 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ed == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_493 <= _ram_T_10;
        end else begin
          ram_493 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_494 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ee == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_494 <= _ram_T_10;
        end else begin
          ram_494 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_495 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ef == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_495 <= _ram_T_10;
        end else begin
          ram_495 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_496 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f0 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_496 <= _ram_T_10;
        end else begin
          ram_496 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_497 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f1 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_497 <= _ram_T_10;
        end else begin
          ram_497 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_498 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f2 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_498 <= _ram_T_10;
        end else begin
          ram_498 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_499 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f3 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_499 <= _ram_T_10;
        end else begin
          ram_499 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_500 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f4 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_500 <= _ram_T_10;
        end else begin
          ram_500 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_501 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f5 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_501 <= _ram_T_10;
        end else begin
          ram_501 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_502 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f6 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_502 <= _ram_T_10;
        end else begin
          ram_502 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_503 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f7 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_503 <= _ram_T_10;
        end else begin
          ram_503 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_504 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f8 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_504 <= _ram_T_10;
        end else begin
          ram_504 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_505 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1f9 == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_505 <= _ram_T_10;
        end else begin
          ram_505 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_506 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1fa == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_506 <= _ram_T_10;
        end else begin
          ram_506 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_507 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1fb == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_507 <= _ram_T_10;
        end else begin
          ram_507 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_508 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1fc == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_508 <= _ram_T_10;
        end else begin
          ram_508 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_509 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1fd == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_509 <= _ram_T_10;
        end else begin
          ram_509 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_510 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1fe == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_510 <= _ram_T_10;
        end else begin
          ram_510 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_511 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (9'h1ff == _GEN_7170) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_511 <= _ram_T_10;
        end else begin
          ram_511 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_512 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h200 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_512 <= _ram_T_10;
        end else begin
          ram_512 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_513 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h201 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_513 <= _ram_T_10;
        end else begin
          ram_513 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_514 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h202 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_514 <= _ram_T_10;
        end else begin
          ram_514 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_515 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h203 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_515 <= _ram_T_10;
        end else begin
          ram_515 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_516 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h204 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_516 <= _ram_T_10;
        end else begin
          ram_516 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_517 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h205 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_517 <= _ram_T_10;
        end else begin
          ram_517 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_518 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h206 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_518 <= _ram_T_10;
        end else begin
          ram_518 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_519 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h207 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_519 <= _ram_T_10;
        end else begin
          ram_519 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_520 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h208 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_520 <= _ram_T_10;
        end else begin
          ram_520 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_521 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h209 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_521 <= _ram_T_10;
        end else begin
          ram_521 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_522 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h20a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_522 <= _ram_T_10;
        end else begin
          ram_522 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_523 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h20b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_523 <= _ram_T_10;
        end else begin
          ram_523 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_524 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h20c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_524 <= _ram_T_10;
        end else begin
          ram_524 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_525 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h20d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_525 <= _ram_T_10;
        end else begin
          ram_525 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_526 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h20e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_526 <= _ram_T_10;
        end else begin
          ram_526 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_527 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h20f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_527 <= _ram_T_10;
        end else begin
          ram_527 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_528 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h210 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_528 <= _ram_T_10;
        end else begin
          ram_528 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_529 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h211 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_529 <= _ram_T_10;
        end else begin
          ram_529 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_530 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h212 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_530 <= _ram_T_10;
        end else begin
          ram_530 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_531 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h213 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_531 <= _ram_T_10;
        end else begin
          ram_531 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_532 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h214 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_532 <= _ram_T_10;
        end else begin
          ram_532 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_533 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h215 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_533 <= _ram_T_10;
        end else begin
          ram_533 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_534 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h216 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_534 <= _ram_T_10;
        end else begin
          ram_534 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_535 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h217 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_535 <= _ram_T_10;
        end else begin
          ram_535 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_536 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h218 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_536 <= _ram_T_10;
        end else begin
          ram_536 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_537 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h219 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_537 <= _ram_T_10;
        end else begin
          ram_537 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_538 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h21a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_538 <= _ram_T_10;
        end else begin
          ram_538 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_539 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h21b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_539 <= _ram_T_10;
        end else begin
          ram_539 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_540 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h21c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_540 <= _ram_T_10;
        end else begin
          ram_540 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_541 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h21d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_541 <= _ram_T_10;
        end else begin
          ram_541 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_542 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h21e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_542 <= _ram_T_10;
        end else begin
          ram_542 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_543 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h21f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_543 <= _ram_T_10;
        end else begin
          ram_543 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_544 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h220 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_544 <= _ram_T_10;
        end else begin
          ram_544 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_545 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h221 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_545 <= _ram_T_10;
        end else begin
          ram_545 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_546 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h222 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_546 <= _ram_T_10;
        end else begin
          ram_546 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_547 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h223 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_547 <= _ram_T_10;
        end else begin
          ram_547 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_548 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h224 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_548 <= _ram_T_10;
        end else begin
          ram_548 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_549 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h225 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_549 <= _ram_T_10;
        end else begin
          ram_549 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_550 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h226 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_550 <= _ram_T_10;
        end else begin
          ram_550 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_551 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h227 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_551 <= _ram_T_10;
        end else begin
          ram_551 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_552 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h228 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_552 <= _ram_T_10;
        end else begin
          ram_552 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_553 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h229 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_553 <= _ram_T_10;
        end else begin
          ram_553 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_554 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h22a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_554 <= _ram_T_10;
        end else begin
          ram_554 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_555 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h22b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_555 <= _ram_T_10;
        end else begin
          ram_555 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_556 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h22c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_556 <= _ram_T_10;
        end else begin
          ram_556 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_557 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h22d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_557 <= _ram_T_10;
        end else begin
          ram_557 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_558 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h22e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_558 <= _ram_T_10;
        end else begin
          ram_558 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_559 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h22f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_559 <= _ram_T_10;
        end else begin
          ram_559 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_560 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h230 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_560 <= _ram_T_10;
        end else begin
          ram_560 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_561 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h231 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_561 <= _ram_T_10;
        end else begin
          ram_561 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_562 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h232 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_562 <= _ram_T_10;
        end else begin
          ram_562 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_563 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h233 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_563 <= _ram_T_10;
        end else begin
          ram_563 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_564 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h234 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_564 <= _ram_T_10;
        end else begin
          ram_564 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_565 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h235 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_565 <= _ram_T_10;
        end else begin
          ram_565 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_566 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h236 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_566 <= _ram_T_10;
        end else begin
          ram_566 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_567 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h237 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_567 <= _ram_T_10;
        end else begin
          ram_567 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_568 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h238 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_568 <= _ram_T_10;
        end else begin
          ram_568 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_569 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h239 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_569 <= _ram_T_10;
        end else begin
          ram_569 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_570 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h23a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_570 <= _ram_T_10;
        end else begin
          ram_570 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_571 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h23b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_571 <= _ram_T_10;
        end else begin
          ram_571 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_572 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h23c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_572 <= _ram_T_10;
        end else begin
          ram_572 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_573 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h23d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_573 <= _ram_T_10;
        end else begin
          ram_573 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_574 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h23e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_574 <= _ram_T_10;
        end else begin
          ram_574 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_575 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h23f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_575 <= _ram_T_10;
        end else begin
          ram_575 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_576 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h240 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_576 <= _ram_T_10;
        end else begin
          ram_576 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_577 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h241 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_577 <= _ram_T_10;
        end else begin
          ram_577 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_578 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h242 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_578 <= _ram_T_10;
        end else begin
          ram_578 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_579 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h243 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_579 <= _ram_T_10;
        end else begin
          ram_579 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_580 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h244 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_580 <= _ram_T_10;
        end else begin
          ram_580 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_581 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h245 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_581 <= _ram_T_10;
        end else begin
          ram_581 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_582 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h246 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_582 <= _ram_T_10;
        end else begin
          ram_582 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_583 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h247 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_583 <= _ram_T_10;
        end else begin
          ram_583 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_584 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h248 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_584 <= _ram_T_10;
        end else begin
          ram_584 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_585 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h249 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_585 <= _ram_T_10;
        end else begin
          ram_585 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_586 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h24a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_586 <= _ram_T_10;
        end else begin
          ram_586 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_587 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h24b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_587 <= _ram_T_10;
        end else begin
          ram_587 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_588 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h24c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_588 <= _ram_T_10;
        end else begin
          ram_588 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_589 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h24d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_589 <= _ram_T_10;
        end else begin
          ram_589 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_590 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h24e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_590 <= _ram_T_10;
        end else begin
          ram_590 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_591 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h24f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_591 <= _ram_T_10;
        end else begin
          ram_591 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_592 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h250 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_592 <= _ram_T_10;
        end else begin
          ram_592 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_593 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h251 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_593 <= _ram_T_10;
        end else begin
          ram_593 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_594 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h252 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_594 <= _ram_T_10;
        end else begin
          ram_594 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_595 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h253 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_595 <= _ram_T_10;
        end else begin
          ram_595 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_596 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h254 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_596 <= _ram_T_10;
        end else begin
          ram_596 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_597 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h255 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_597 <= _ram_T_10;
        end else begin
          ram_597 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_598 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h256 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_598 <= _ram_T_10;
        end else begin
          ram_598 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_599 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h257 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_599 <= _ram_T_10;
        end else begin
          ram_599 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_600 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h258 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_600 <= _ram_T_10;
        end else begin
          ram_600 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_601 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h259 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_601 <= _ram_T_10;
        end else begin
          ram_601 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_602 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h25a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_602 <= _ram_T_10;
        end else begin
          ram_602 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_603 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h25b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_603 <= _ram_T_10;
        end else begin
          ram_603 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_604 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h25c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_604 <= _ram_T_10;
        end else begin
          ram_604 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_605 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h25d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_605 <= _ram_T_10;
        end else begin
          ram_605 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_606 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h25e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_606 <= _ram_T_10;
        end else begin
          ram_606 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_607 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h25f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_607 <= _ram_T_10;
        end else begin
          ram_607 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_608 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h260 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_608 <= _ram_T_10;
        end else begin
          ram_608 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_609 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h261 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_609 <= _ram_T_10;
        end else begin
          ram_609 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_610 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h262 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_610 <= _ram_T_10;
        end else begin
          ram_610 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_611 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h263 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_611 <= _ram_T_10;
        end else begin
          ram_611 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_612 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h264 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_612 <= _ram_T_10;
        end else begin
          ram_612 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_613 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h265 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_613 <= _ram_T_10;
        end else begin
          ram_613 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_614 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h266 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_614 <= _ram_T_10;
        end else begin
          ram_614 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_615 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h267 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_615 <= _ram_T_10;
        end else begin
          ram_615 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_616 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h268 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_616 <= _ram_T_10;
        end else begin
          ram_616 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_617 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h269 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_617 <= _ram_T_10;
        end else begin
          ram_617 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_618 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h26a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_618 <= _ram_T_10;
        end else begin
          ram_618 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_619 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h26b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_619 <= _ram_T_10;
        end else begin
          ram_619 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_620 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h26c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_620 <= _ram_T_10;
        end else begin
          ram_620 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_621 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h26d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_621 <= _ram_T_10;
        end else begin
          ram_621 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_622 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h26e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_622 <= _ram_T_10;
        end else begin
          ram_622 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_623 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h26f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_623 <= _ram_T_10;
        end else begin
          ram_623 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_624 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h270 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_624 <= _ram_T_10;
        end else begin
          ram_624 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_625 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h271 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_625 <= _ram_T_10;
        end else begin
          ram_625 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_626 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h272 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_626 <= _ram_T_10;
        end else begin
          ram_626 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_627 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h273 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_627 <= _ram_T_10;
        end else begin
          ram_627 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_628 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h274 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_628 <= _ram_T_10;
        end else begin
          ram_628 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_629 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h275 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_629 <= _ram_T_10;
        end else begin
          ram_629 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_630 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h276 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_630 <= _ram_T_10;
        end else begin
          ram_630 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_631 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h277 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_631 <= _ram_T_10;
        end else begin
          ram_631 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_632 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h278 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_632 <= _ram_T_10;
        end else begin
          ram_632 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_633 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h279 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_633 <= _ram_T_10;
        end else begin
          ram_633 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_634 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h27a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_634 <= _ram_T_10;
        end else begin
          ram_634 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_635 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h27b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_635 <= _ram_T_10;
        end else begin
          ram_635 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_636 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h27c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_636 <= _ram_T_10;
        end else begin
          ram_636 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_637 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h27d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_637 <= _ram_T_10;
        end else begin
          ram_637 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_638 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h27e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_638 <= _ram_T_10;
        end else begin
          ram_638 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_639 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h27f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_639 <= _ram_T_10;
        end else begin
          ram_639 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_640 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h280 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_640 <= _ram_T_10;
        end else begin
          ram_640 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_641 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h281 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_641 <= _ram_T_10;
        end else begin
          ram_641 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_642 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h282 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_642 <= _ram_T_10;
        end else begin
          ram_642 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_643 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h283 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_643 <= _ram_T_10;
        end else begin
          ram_643 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_644 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h284 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_644 <= _ram_T_10;
        end else begin
          ram_644 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_645 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h285 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_645 <= _ram_T_10;
        end else begin
          ram_645 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_646 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h286 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_646 <= _ram_T_10;
        end else begin
          ram_646 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_647 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h287 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_647 <= _ram_T_10;
        end else begin
          ram_647 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_648 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h288 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_648 <= _ram_T_10;
        end else begin
          ram_648 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_649 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h289 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_649 <= _ram_T_10;
        end else begin
          ram_649 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_650 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h28a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_650 <= _ram_T_10;
        end else begin
          ram_650 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_651 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h28b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_651 <= _ram_T_10;
        end else begin
          ram_651 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_652 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h28c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_652 <= _ram_T_10;
        end else begin
          ram_652 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_653 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h28d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_653 <= _ram_T_10;
        end else begin
          ram_653 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_654 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h28e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_654 <= _ram_T_10;
        end else begin
          ram_654 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_655 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h28f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_655 <= _ram_T_10;
        end else begin
          ram_655 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_656 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h290 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_656 <= _ram_T_10;
        end else begin
          ram_656 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_657 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h291 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_657 <= _ram_T_10;
        end else begin
          ram_657 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_658 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h292 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_658 <= _ram_T_10;
        end else begin
          ram_658 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_659 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h293 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_659 <= _ram_T_10;
        end else begin
          ram_659 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_660 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h294 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_660 <= _ram_T_10;
        end else begin
          ram_660 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_661 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h295 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_661 <= _ram_T_10;
        end else begin
          ram_661 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_662 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h296 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_662 <= _ram_T_10;
        end else begin
          ram_662 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_663 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h297 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_663 <= _ram_T_10;
        end else begin
          ram_663 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_664 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h298 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_664 <= _ram_T_10;
        end else begin
          ram_664 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_665 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h299 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_665 <= _ram_T_10;
        end else begin
          ram_665 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_666 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h29a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_666 <= _ram_T_10;
        end else begin
          ram_666 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_667 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h29b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_667 <= _ram_T_10;
        end else begin
          ram_667 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_668 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h29c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_668 <= _ram_T_10;
        end else begin
          ram_668 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_669 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h29d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_669 <= _ram_T_10;
        end else begin
          ram_669 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_670 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h29e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_670 <= _ram_T_10;
        end else begin
          ram_670 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_671 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h29f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_671 <= _ram_T_10;
        end else begin
          ram_671 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_672 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_672 <= _ram_T_10;
        end else begin
          ram_672 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_673 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_673 <= _ram_T_10;
        end else begin
          ram_673 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_674 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_674 <= _ram_T_10;
        end else begin
          ram_674 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_675 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_675 <= _ram_T_10;
        end else begin
          ram_675 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_676 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_676 <= _ram_T_10;
        end else begin
          ram_676 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_677 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_677 <= _ram_T_10;
        end else begin
          ram_677 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_678 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_678 <= _ram_T_10;
        end else begin
          ram_678 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_679 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_679 <= _ram_T_10;
        end else begin
          ram_679 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_680 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_680 <= _ram_T_10;
        end else begin
          ram_680 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_681 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2a9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_681 <= _ram_T_10;
        end else begin
          ram_681 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_682 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2aa == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_682 <= _ram_T_10;
        end else begin
          ram_682 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_683 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ab == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_683 <= _ram_T_10;
        end else begin
          ram_683 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_684 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ac == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_684 <= _ram_T_10;
        end else begin
          ram_684 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_685 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ad == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_685 <= _ram_T_10;
        end else begin
          ram_685 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_686 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ae == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_686 <= _ram_T_10;
        end else begin
          ram_686 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_687 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2af == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_687 <= _ram_T_10;
        end else begin
          ram_687 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_688 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_688 <= _ram_T_10;
        end else begin
          ram_688 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_689 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_689 <= _ram_T_10;
        end else begin
          ram_689 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_690 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_690 <= _ram_T_10;
        end else begin
          ram_690 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_691 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_691 <= _ram_T_10;
        end else begin
          ram_691 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_692 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_692 <= _ram_T_10;
        end else begin
          ram_692 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_693 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_693 <= _ram_T_10;
        end else begin
          ram_693 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_694 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_694 <= _ram_T_10;
        end else begin
          ram_694 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_695 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_695 <= _ram_T_10;
        end else begin
          ram_695 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_696 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_696 <= _ram_T_10;
        end else begin
          ram_696 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_697 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2b9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_697 <= _ram_T_10;
        end else begin
          ram_697 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_698 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ba == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_698 <= _ram_T_10;
        end else begin
          ram_698 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_699 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2bb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_699 <= _ram_T_10;
        end else begin
          ram_699 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_700 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2bc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_700 <= _ram_T_10;
        end else begin
          ram_700 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_701 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2bd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_701 <= _ram_T_10;
        end else begin
          ram_701 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_702 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2be == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_702 <= _ram_T_10;
        end else begin
          ram_702 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_703 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2bf == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_703 <= _ram_T_10;
        end else begin
          ram_703 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_704 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_704 <= _ram_T_10;
        end else begin
          ram_704 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_705 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_705 <= _ram_T_10;
        end else begin
          ram_705 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_706 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_706 <= _ram_T_10;
        end else begin
          ram_706 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_707 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_707 <= _ram_T_10;
        end else begin
          ram_707 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_708 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_708 <= _ram_T_10;
        end else begin
          ram_708 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_709 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_709 <= _ram_T_10;
        end else begin
          ram_709 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_710 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_710 <= _ram_T_10;
        end else begin
          ram_710 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_711 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_711 <= _ram_T_10;
        end else begin
          ram_711 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_712 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_712 <= _ram_T_10;
        end else begin
          ram_712 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_713 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2c9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_713 <= _ram_T_10;
        end else begin
          ram_713 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_714 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ca == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_714 <= _ram_T_10;
        end else begin
          ram_714 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_715 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2cb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_715 <= _ram_T_10;
        end else begin
          ram_715 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_716 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2cc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_716 <= _ram_T_10;
        end else begin
          ram_716 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_717 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2cd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_717 <= _ram_T_10;
        end else begin
          ram_717 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_718 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ce == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_718 <= _ram_T_10;
        end else begin
          ram_718 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_719 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2cf == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_719 <= _ram_T_10;
        end else begin
          ram_719 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_720 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_720 <= _ram_T_10;
        end else begin
          ram_720 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_721 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_721 <= _ram_T_10;
        end else begin
          ram_721 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_722 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_722 <= _ram_T_10;
        end else begin
          ram_722 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_723 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_723 <= _ram_T_10;
        end else begin
          ram_723 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_724 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_724 <= _ram_T_10;
        end else begin
          ram_724 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_725 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_725 <= _ram_T_10;
        end else begin
          ram_725 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_726 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_726 <= _ram_T_10;
        end else begin
          ram_726 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_727 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_727 <= _ram_T_10;
        end else begin
          ram_727 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_728 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_728 <= _ram_T_10;
        end else begin
          ram_728 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_729 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2d9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_729 <= _ram_T_10;
        end else begin
          ram_729 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_730 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2da == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_730 <= _ram_T_10;
        end else begin
          ram_730 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_731 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2db == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_731 <= _ram_T_10;
        end else begin
          ram_731 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_732 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2dc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_732 <= _ram_T_10;
        end else begin
          ram_732 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_733 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2dd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_733 <= _ram_T_10;
        end else begin
          ram_733 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_734 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2de == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_734 <= _ram_T_10;
        end else begin
          ram_734 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_735 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2df == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_735 <= _ram_T_10;
        end else begin
          ram_735 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_736 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_736 <= _ram_T_10;
        end else begin
          ram_736 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_737 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_737 <= _ram_T_10;
        end else begin
          ram_737 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_738 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_738 <= _ram_T_10;
        end else begin
          ram_738 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_739 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_739 <= _ram_T_10;
        end else begin
          ram_739 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_740 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_740 <= _ram_T_10;
        end else begin
          ram_740 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_741 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_741 <= _ram_T_10;
        end else begin
          ram_741 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_742 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_742 <= _ram_T_10;
        end else begin
          ram_742 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_743 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_743 <= _ram_T_10;
        end else begin
          ram_743 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_744 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_744 <= _ram_T_10;
        end else begin
          ram_744 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_745 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2e9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_745 <= _ram_T_10;
        end else begin
          ram_745 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_746 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ea == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_746 <= _ram_T_10;
        end else begin
          ram_746 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_747 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2eb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_747 <= _ram_T_10;
        end else begin
          ram_747 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_748 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ec == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_748 <= _ram_T_10;
        end else begin
          ram_748 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_749 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ed == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_749 <= _ram_T_10;
        end else begin
          ram_749 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_750 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ee == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_750 <= _ram_T_10;
        end else begin
          ram_750 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_751 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ef == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_751 <= _ram_T_10;
        end else begin
          ram_751 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_752 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_752 <= _ram_T_10;
        end else begin
          ram_752 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_753 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_753 <= _ram_T_10;
        end else begin
          ram_753 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_754 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_754 <= _ram_T_10;
        end else begin
          ram_754 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_755 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_755 <= _ram_T_10;
        end else begin
          ram_755 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_756 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_756 <= _ram_T_10;
        end else begin
          ram_756 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_757 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_757 <= _ram_T_10;
        end else begin
          ram_757 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_758 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_758 <= _ram_T_10;
        end else begin
          ram_758 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_759 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_759 <= _ram_T_10;
        end else begin
          ram_759 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_760 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_760 <= _ram_T_10;
        end else begin
          ram_760 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_761 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2f9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_761 <= _ram_T_10;
        end else begin
          ram_761 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_762 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2fa == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_762 <= _ram_T_10;
        end else begin
          ram_762 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_763 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2fb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_763 <= _ram_T_10;
        end else begin
          ram_763 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_764 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2fc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_764 <= _ram_T_10;
        end else begin
          ram_764 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_765 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2fd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_765 <= _ram_T_10;
        end else begin
          ram_765 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_766 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2fe == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_766 <= _ram_T_10;
        end else begin
          ram_766 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_767 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h2ff == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_767 <= _ram_T_10;
        end else begin
          ram_767 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_768 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h300 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_768 <= _ram_T_10;
        end else begin
          ram_768 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_769 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h301 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_769 <= _ram_T_10;
        end else begin
          ram_769 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_770 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h302 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_770 <= _ram_T_10;
        end else begin
          ram_770 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_771 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h303 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_771 <= _ram_T_10;
        end else begin
          ram_771 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_772 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h304 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_772 <= _ram_T_10;
        end else begin
          ram_772 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_773 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h305 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_773 <= _ram_T_10;
        end else begin
          ram_773 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_774 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h306 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_774 <= _ram_T_10;
        end else begin
          ram_774 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_775 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h307 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_775 <= _ram_T_10;
        end else begin
          ram_775 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_776 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h308 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_776 <= _ram_T_10;
        end else begin
          ram_776 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_777 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h309 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_777 <= _ram_T_10;
        end else begin
          ram_777 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_778 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h30a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_778 <= _ram_T_10;
        end else begin
          ram_778 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_779 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h30b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_779 <= _ram_T_10;
        end else begin
          ram_779 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_780 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h30c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_780 <= _ram_T_10;
        end else begin
          ram_780 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_781 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h30d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_781 <= _ram_T_10;
        end else begin
          ram_781 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_782 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h30e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_782 <= _ram_T_10;
        end else begin
          ram_782 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_783 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h30f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_783 <= _ram_T_10;
        end else begin
          ram_783 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_784 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h310 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_784 <= _ram_T_10;
        end else begin
          ram_784 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_785 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h311 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_785 <= _ram_T_10;
        end else begin
          ram_785 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_786 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h312 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_786 <= _ram_T_10;
        end else begin
          ram_786 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_787 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h313 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_787 <= _ram_T_10;
        end else begin
          ram_787 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_788 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h314 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_788 <= _ram_T_10;
        end else begin
          ram_788 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_789 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h315 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_789 <= _ram_T_10;
        end else begin
          ram_789 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_790 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h316 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_790 <= _ram_T_10;
        end else begin
          ram_790 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_791 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h317 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_791 <= _ram_T_10;
        end else begin
          ram_791 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_792 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h318 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_792 <= _ram_T_10;
        end else begin
          ram_792 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_793 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h319 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_793 <= _ram_T_10;
        end else begin
          ram_793 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_794 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h31a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_794 <= _ram_T_10;
        end else begin
          ram_794 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_795 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h31b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_795 <= _ram_T_10;
        end else begin
          ram_795 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_796 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h31c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_796 <= _ram_T_10;
        end else begin
          ram_796 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_797 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h31d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_797 <= _ram_T_10;
        end else begin
          ram_797 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_798 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h31e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_798 <= _ram_T_10;
        end else begin
          ram_798 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_799 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h31f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_799 <= _ram_T_10;
        end else begin
          ram_799 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_800 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h320 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_800 <= _ram_T_10;
        end else begin
          ram_800 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_801 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h321 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_801 <= _ram_T_10;
        end else begin
          ram_801 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_802 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h322 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_802 <= _ram_T_10;
        end else begin
          ram_802 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_803 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h323 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_803 <= _ram_T_10;
        end else begin
          ram_803 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_804 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h324 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_804 <= _ram_T_10;
        end else begin
          ram_804 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_805 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h325 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_805 <= _ram_T_10;
        end else begin
          ram_805 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_806 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h326 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_806 <= _ram_T_10;
        end else begin
          ram_806 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_807 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h327 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_807 <= _ram_T_10;
        end else begin
          ram_807 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_808 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h328 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_808 <= _ram_T_10;
        end else begin
          ram_808 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_809 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h329 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_809 <= _ram_T_10;
        end else begin
          ram_809 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_810 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h32a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_810 <= _ram_T_10;
        end else begin
          ram_810 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_811 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h32b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_811 <= _ram_T_10;
        end else begin
          ram_811 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_812 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h32c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_812 <= _ram_T_10;
        end else begin
          ram_812 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_813 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h32d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_813 <= _ram_T_10;
        end else begin
          ram_813 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_814 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h32e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_814 <= _ram_T_10;
        end else begin
          ram_814 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_815 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h32f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_815 <= _ram_T_10;
        end else begin
          ram_815 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_816 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h330 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_816 <= _ram_T_10;
        end else begin
          ram_816 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_817 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h331 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_817 <= _ram_T_10;
        end else begin
          ram_817 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_818 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h332 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_818 <= _ram_T_10;
        end else begin
          ram_818 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_819 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h333 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_819 <= _ram_T_10;
        end else begin
          ram_819 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_820 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h334 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_820 <= _ram_T_10;
        end else begin
          ram_820 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_821 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h335 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_821 <= _ram_T_10;
        end else begin
          ram_821 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_822 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h336 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_822 <= _ram_T_10;
        end else begin
          ram_822 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_823 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h337 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_823 <= _ram_T_10;
        end else begin
          ram_823 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_824 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h338 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_824 <= _ram_T_10;
        end else begin
          ram_824 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_825 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h339 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_825 <= _ram_T_10;
        end else begin
          ram_825 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_826 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h33a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_826 <= _ram_T_10;
        end else begin
          ram_826 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_827 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h33b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_827 <= _ram_T_10;
        end else begin
          ram_827 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_828 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h33c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_828 <= _ram_T_10;
        end else begin
          ram_828 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_829 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h33d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_829 <= _ram_T_10;
        end else begin
          ram_829 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_830 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h33e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_830 <= _ram_T_10;
        end else begin
          ram_830 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_831 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h33f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_831 <= _ram_T_10;
        end else begin
          ram_831 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_832 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h340 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_832 <= _ram_T_10;
        end else begin
          ram_832 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_833 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h341 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_833 <= _ram_T_10;
        end else begin
          ram_833 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_834 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h342 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_834 <= _ram_T_10;
        end else begin
          ram_834 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_835 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h343 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_835 <= _ram_T_10;
        end else begin
          ram_835 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_836 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h344 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_836 <= _ram_T_10;
        end else begin
          ram_836 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_837 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h345 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_837 <= _ram_T_10;
        end else begin
          ram_837 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_838 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h346 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_838 <= _ram_T_10;
        end else begin
          ram_838 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_839 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h347 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_839 <= _ram_T_10;
        end else begin
          ram_839 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_840 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h348 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_840 <= _ram_T_10;
        end else begin
          ram_840 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_841 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h349 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_841 <= _ram_T_10;
        end else begin
          ram_841 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_842 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h34a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_842 <= _ram_T_10;
        end else begin
          ram_842 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_843 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h34b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_843 <= _ram_T_10;
        end else begin
          ram_843 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_844 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h34c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_844 <= _ram_T_10;
        end else begin
          ram_844 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_845 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h34d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_845 <= _ram_T_10;
        end else begin
          ram_845 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_846 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h34e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_846 <= _ram_T_10;
        end else begin
          ram_846 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_847 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h34f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_847 <= _ram_T_10;
        end else begin
          ram_847 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_848 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h350 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_848 <= _ram_T_10;
        end else begin
          ram_848 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_849 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h351 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_849 <= _ram_T_10;
        end else begin
          ram_849 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_850 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h352 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_850 <= _ram_T_10;
        end else begin
          ram_850 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_851 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h353 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_851 <= _ram_T_10;
        end else begin
          ram_851 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_852 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h354 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_852 <= _ram_T_10;
        end else begin
          ram_852 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_853 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h355 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_853 <= _ram_T_10;
        end else begin
          ram_853 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_854 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h356 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_854 <= _ram_T_10;
        end else begin
          ram_854 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_855 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h357 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_855 <= _ram_T_10;
        end else begin
          ram_855 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_856 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h358 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_856 <= _ram_T_10;
        end else begin
          ram_856 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_857 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h359 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_857 <= _ram_T_10;
        end else begin
          ram_857 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_858 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h35a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_858 <= _ram_T_10;
        end else begin
          ram_858 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_859 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h35b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_859 <= _ram_T_10;
        end else begin
          ram_859 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_860 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h35c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_860 <= _ram_T_10;
        end else begin
          ram_860 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_861 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h35d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_861 <= _ram_T_10;
        end else begin
          ram_861 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_862 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h35e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_862 <= _ram_T_10;
        end else begin
          ram_862 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_863 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h35f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_863 <= _ram_T_10;
        end else begin
          ram_863 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_864 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h360 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_864 <= _ram_T_10;
        end else begin
          ram_864 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_865 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h361 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_865 <= _ram_T_10;
        end else begin
          ram_865 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_866 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h362 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_866 <= _ram_T_10;
        end else begin
          ram_866 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_867 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h363 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_867 <= _ram_T_10;
        end else begin
          ram_867 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_868 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h364 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_868 <= _ram_T_10;
        end else begin
          ram_868 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_869 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h365 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_869 <= _ram_T_10;
        end else begin
          ram_869 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_870 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h366 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_870 <= _ram_T_10;
        end else begin
          ram_870 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_871 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h367 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_871 <= _ram_T_10;
        end else begin
          ram_871 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_872 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h368 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_872 <= _ram_T_10;
        end else begin
          ram_872 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_873 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h369 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_873 <= _ram_T_10;
        end else begin
          ram_873 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_874 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h36a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_874 <= _ram_T_10;
        end else begin
          ram_874 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_875 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h36b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_875 <= _ram_T_10;
        end else begin
          ram_875 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_876 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h36c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_876 <= _ram_T_10;
        end else begin
          ram_876 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_877 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h36d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_877 <= _ram_T_10;
        end else begin
          ram_877 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_878 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h36e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_878 <= _ram_T_10;
        end else begin
          ram_878 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_879 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h36f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_879 <= _ram_T_10;
        end else begin
          ram_879 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_880 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h370 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_880 <= _ram_T_10;
        end else begin
          ram_880 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_881 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h371 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_881 <= _ram_T_10;
        end else begin
          ram_881 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_882 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h372 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_882 <= _ram_T_10;
        end else begin
          ram_882 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_883 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h373 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_883 <= _ram_T_10;
        end else begin
          ram_883 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_884 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h374 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_884 <= _ram_T_10;
        end else begin
          ram_884 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_885 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h375 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_885 <= _ram_T_10;
        end else begin
          ram_885 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_886 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h376 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_886 <= _ram_T_10;
        end else begin
          ram_886 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_887 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h377 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_887 <= _ram_T_10;
        end else begin
          ram_887 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_888 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h378 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_888 <= _ram_T_10;
        end else begin
          ram_888 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_889 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h379 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_889 <= _ram_T_10;
        end else begin
          ram_889 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_890 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h37a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_890 <= _ram_T_10;
        end else begin
          ram_890 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_891 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h37b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_891 <= _ram_T_10;
        end else begin
          ram_891 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_892 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h37c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_892 <= _ram_T_10;
        end else begin
          ram_892 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_893 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h37d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_893 <= _ram_T_10;
        end else begin
          ram_893 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_894 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h37e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_894 <= _ram_T_10;
        end else begin
          ram_894 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_895 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h37f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_895 <= _ram_T_10;
        end else begin
          ram_895 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_896 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h380 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_896 <= _ram_T_10;
        end else begin
          ram_896 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_897 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h381 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_897 <= _ram_T_10;
        end else begin
          ram_897 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_898 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h382 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_898 <= _ram_T_10;
        end else begin
          ram_898 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_899 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h383 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_899 <= _ram_T_10;
        end else begin
          ram_899 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_900 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h384 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_900 <= _ram_T_10;
        end else begin
          ram_900 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_901 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h385 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_901 <= _ram_T_10;
        end else begin
          ram_901 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_902 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h386 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_902 <= _ram_T_10;
        end else begin
          ram_902 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_903 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h387 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_903 <= _ram_T_10;
        end else begin
          ram_903 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_904 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h388 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_904 <= _ram_T_10;
        end else begin
          ram_904 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_905 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h389 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_905 <= _ram_T_10;
        end else begin
          ram_905 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_906 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h38a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_906 <= _ram_T_10;
        end else begin
          ram_906 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_907 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h38b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_907 <= _ram_T_10;
        end else begin
          ram_907 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_908 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h38c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_908 <= _ram_T_10;
        end else begin
          ram_908 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_909 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h38d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_909 <= _ram_T_10;
        end else begin
          ram_909 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_910 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h38e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_910 <= _ram_T_10;
        end else begin
          ram_910 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_911 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h38f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_911 <= _ram_T_10;
        end else begin
          ram_911 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_912 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h390 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_912 <= _ram_T_10;
        end else begin
          ram_912 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_913 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h391 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_913 <= _ram_T_10;
        end else begin
          ram_913 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_914 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h392 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_914 <= _ram_T_10;
        end else begin
          ram_914 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_915 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h393 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_915 <= _ram_T_10;
        end else begin
          ram_915 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_916 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h394 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_916 <= _ram_T_10;
        end else begin
          ram_916 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_917 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h395 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_917 <= _ram_T_10;
        end else begin
          ram_917 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_918 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h396 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_918 <= _ram_T_10;
        end else begin
          ram_918 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_919 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h397 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_919 <= _ram_T_10;
        end else begin
          ram_919 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_920 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h398 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_920 <= _ram_T_10;
        end else begin
          ram_920 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_921 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h399 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_921 <= _ram_T_10;
        end else begin
          ram_921 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_922 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h39a == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_922 <= _ram_T_10;
        end else begin
          ram_922 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_923 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h39b == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_923 <= _ram_T_10;
        end else begin
          ram_923 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_924 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h39c == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_924 <= _ram_T_10;
        end else begin
          ram_924 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_925 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h39d == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_925 <= _ram_T_10;
        end else begin
          ram_925 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_926 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h39e == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_926 <= _ram_T_10;
        end else begin
          ram_926 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_927 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h39f == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_927 <= _ram_T_10;
        end else begin
          ram_927 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_928 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_928 <= _ram_T_10;
        end else begin
          ram_928 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_929 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_929 <= _ram_T_10;
        end else begin
          ram_929 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_930 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_930 <= _ram_T_10;
        end else begin
          ram_930 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_931 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_931 <= _ram_T_10;
        end else begin
          ram_931 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_932 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_932 <= _ram_T_10;
        end else begin
          ram_932 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_933 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_933 <= _ram_T_10;
        end else begin
          ram_933 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_934 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_934 <= _ram_T_10;
        end else begin
          ram_934 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_935 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_935 <= _ram_T_10;
        end else begin
          ram_935 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_936 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_936 <= _ram_T_10;
        end else begin
          ram_936 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_937 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3a9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_937 <= _ram_T_10;
        end else begin
          ram_937 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_938 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3aa == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_938 <= _ram_T_10;
        end else begin
          ram_938 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_939 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ab == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_939 <= _ram_T_10;
        end else begin
          ram_939 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_940 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ac == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_940 <= _ram_T_10;
        end else begin
          ram_940 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_941 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ad == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_941 <= _ram_T_10;
        end else begin
          ram_941 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_942 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ae == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_942 <= _ram_T_10;
        end else begin
          ram_942 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_943 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3af == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_943 <= _ram_T_10;
        end else begin
          ram_943 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_944 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_944 <= _ram_T_10;
        end else begin
          ram_944 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_945 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_945 <= _ram_T_10;
        end else begin
          ram_945 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_946 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_946 <= _ram_T_10;
        end else begin
          ram_946 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_947 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_947 <= _ram_T_10;
        end else begin
          ram_947 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_948 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_948 <= _ram_T_10;
        end else begin
          ram_948 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_949 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_949 <= _ram_T_10;
        end else begin
          ram_949 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_950 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_950 <= _ram_T_10;
        end else begin
          ram_950 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_951 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_951 <= _ram_T_10;
        end else begin
          ram_951 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_952 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_952 <= _ram_T_10;
        end else begin
          ram_952 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_953 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3b9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_953 <= _ram_T_10;
        end else begin
          ram_953 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_954 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ba == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_954 <= _ram_T_10;
        end else begin
          ram_954 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_955 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3bb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_955 <= _ram_T_10;
        end else begin
          ram_955 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_956 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3bc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_956 <= _ram_T_10;
        end else begin
          ram_956 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_957 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3bd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_957 <= _ram_T_10;
        end else begin
          ram_957 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_958 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3be == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_958 <= _ram_T_10;
        end else begin
          ram_958 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_959 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3bf == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_959 <= _ram_T_10;
        end else begin
          ram_959 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_960 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_960 <= _ram_T_10;
        end else begin
          ram_960 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_961 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_961 <= _ram_T_10;
        end else begin
          ram_961 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_962 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_962 <= _ram_T_10;
        end else begin
          ram_962 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_963 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_963 <= _ram_T_10;
        end else begin
          ram_963 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_964 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_964 <= _ram_T_10;
        end else begin
          ram_964 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_965 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_965 <= _ram_T_10;
        end else begin
          ram_965 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_966 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_966 <= _ram_T_10;
        end else begin
          ram_966 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_967 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_967 <= _ram_T_10;
        end else begin
          ram_967 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_968 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_968 <= _ram_T_10;
        end else begin
          ram_968 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_969 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3c9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_969 <= _ram_T_10;
        end else begin
          ram_969 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_970 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ca == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_970 <= _ram_T_10;
        end else begin
          ram_970 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_971 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3cb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_971 <= _ram_T_10;
        end else begin
          ram_971 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_972 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3cc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_972 <= _ram_T_10;
        end else begin
          ram_972 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_973 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3cd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_973 <= _ram_T_10;
        end else begin
          ram_973 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_974 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ce == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_974 <= _ram_T_10;
        end else begin
          ram_974 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_975 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3cf == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_975 <= _ram_T_10;
        end else begin
          ram_975 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_976 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_976 <= _ram_T_10;
        end else begin
          ram_976 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_977 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_977 <= _ram_T_10;
        end else begin
          ram_977 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_978 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_978 <= _ram_T_10;
        end else begin
          ram_978 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_979 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_979 <= _ram_T_10;
        end else begin
          ram_979 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_980 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_980 <= _ram_T_10;
        end else begin
          ram_980 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_981 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_981 <= _ram_T_10;
        end else begin
          ram_981 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_982 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_982 <= _ram_T_10;
        end else begin
          ram_982 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_983 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_983 <= _ram_T_10;
        end else begin
          ram_983 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_984 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_984 <= _ram_T_10;
        end else begin
          ram_984 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_985 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3d9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_985 <= _ram_T_10;
        end else begin
          ram_985 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_986 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3da == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_986 <= _ram_T_10;
        end else begin
          ram_986 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_987 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3db == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_987 <= _ram_T_10;
        end else begin
          ram_987 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_988 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3dc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_988 <= _ram_T_10;
        end else begin
          ram_988 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_989 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3dd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_989 <= _ram_T_10;
        end else begin
          ram_989 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_990 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3de == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_990 <= _ram_T_10;
        end else begin
          ram_990 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_991 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3df == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_991 <= _ram_T_10;
        end else begin
          ram_991 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_992 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_992 <= _ram_T_10;
        end else begin
          ram_992 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_993 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_993 <= _ram_T_10;
        end else begin
          ram_993 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_994 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_994 <= _ram_T_10;
        end else begin
          ram_994 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_995 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_995 <= _ram_T_10;
        end else begin
          ram_995 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_996 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_996 <= _ram_T_10;
        end else begin
          ram_996 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_997 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_997 <= _ram_T_10;
        end else begin
          ram_997 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_998 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_998 <= _ram_T_10;
        end else begin
          ram_998 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_999 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_999 <= _ram_T_10;
        end else begin
          ram_999 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1000 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1000 <= _ram_T_10;
        end else begin
          ram_1000 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1001 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3e9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1001 <= _ram_T_10;
        end else begin
          ram_1001 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1002 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ea == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1002 <= _ram_T_10;
        end else begin
          ram_1002 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1003 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3eb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1003 <= _ram_T_10;
        end else begin
          ram_1003 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1004 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ec == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1004 <= _ram_T_10;
        end else begin
          ram_1004 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1005 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ed == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1005 <= _ram_T_10;
        end else begin
          ram_1005 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1006 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ee == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1006 <= _ram_T_10;
        end else begin
          ram_1006 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1007 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ef == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1007 <= _ram_T_10;
        end else begin
          ram_1007 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1008 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f0 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1008 <= _ram_T_10;
        end else begin
          ram_1008 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1009 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f1 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1009 <= _ram_T_10;
        end else begin
          ram_1009 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1010 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f2 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1010 <= _ram_T_10;
        end else begin
          ram_1010 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1011 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f3 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1011 <= _ram_T_10;
        end else begin
          ram_1011 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1012 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f4 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1012 <= _ram_T_10;
        end else begin
          ram_1012 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1013 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f5 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1013 <= _ram_T_10;
        end else begin
          ram_1013 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1014 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f6 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1014 <= _ram_T_10;
        end else begin
          ram_1014 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1015 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f7 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1015 <= _ram_T_10;
        end else begin
          ram_1015 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1016 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f8 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1016 <= _ram_T_10;
        end else begin
          ram_1016 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1017 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3f9 == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1017 <= _ram_T_10;
        end else begin
          ram_1017 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1018 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3fa == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1018 <= _ram_T_10;
        end else begin
          ram_1018 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1019 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3fb == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1019 <= _ram_T_10;
        end else begin
          ram_1019 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1020 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3fc == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1020 <= _ram_T_10;
        end else begin
          ram_1020 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1021 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3fd == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1021 <= _ram_T_10;
        end else begin
          ram_1021 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1022 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3fe == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1022 <= _ram_T_10;
        end else begin
          ram_1022 <= _ram_T_14;
        end
      end
    end
    if (reset) begin // @[DataMemory.scala 26:20]
      ram_1023 <= 32'h0; // @[DataMemory.scala 26:20]
    end else if (io_writeEnable) begin // @[DataMemory.scala 64:24]
      if (10'h3ff == _GEN_7426) begin // @[DataMemory.scala 67:18]
        if (2'h3 == io_addr[1:0]) begin // @[Mux.scala 81:58]
          ram_1023 <= _ram_T_10;
        end else begin
          ram_1023 <= _ram_T_14;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ram_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ram_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  ram_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  ram_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  ram_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  ram_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  ram_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ram_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  ram_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  ram_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  ram_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  ram_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  ram_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  ram_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  ram_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  ram_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  ram_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  ram_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  ram_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  ram_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  ram_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  ram_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  ram_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  ram_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  ram_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  ram_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  ram_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  ram_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  ram_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  ram_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  ram_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  ram_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  ram_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  ram_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  ram_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  ram_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  ram_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  ram_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  ram_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  ram_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  ram_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  ram_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  ram_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  ram_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  ram_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  ram_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  ram_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  ram_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  ram_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  ram_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  ram_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  ram_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  ram_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  ram_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  ram_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  ram_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  ram_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  ram_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  ram_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  ram_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  ram_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  ram_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  ram_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  ram_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  ram_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  ram_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  ram_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  ram_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  ram_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  ram_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  ram_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  ram_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  ram_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  ram_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  ram_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  ram_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  ram_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  ram_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  ram_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  ram_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  ram_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  ram_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  ram_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  ram_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  ram_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  ram_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  ram_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  ram_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  ram_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  ram_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  ram_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  ram_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  ram_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  ram_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  ram_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  ram_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  ram_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  ram_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  ram_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  ram_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  ram_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  ram_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  ram_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  ram_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  ram_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  ram_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  ram_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  ram_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  ram_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  ram_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  ram_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  ram_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  ram_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  ram_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  ram_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  ram_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  ram_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  ram_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  ram_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  ram_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  ram_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  ram_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  ram_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  ram_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  ram_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  ram_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  ram_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  ram_127 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  ram_128 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  ram_129 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  ram_130 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  ram_131 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  ram_132 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  ram_133 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  ram_134 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  ram_135 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  ram_136 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  ram_137 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  ram_138 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  ram_139 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  ram_140 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  ram_141 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  ram_142 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  ram_143 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  ram_144 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  ram_145 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  ram_146 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  ram_147 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  ram_148 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  ram_149 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  ram_150 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  ram_151 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  ram_152 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  ram_153 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  ram_154 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  ram_155 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  ram_156 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  ram_157 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  ram_158 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  ram_159 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  ram_160 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  ram_161 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  ram_162 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  ram_163 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  ram_164 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ram_165 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ram_166 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ram_167 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ram_168 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ram_169 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ram_170 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ram_171 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ram_172 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ram_173 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ram_174 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ram_175 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ram_176 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ram_177 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ram_178 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ram_179 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ram_180 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ram_181 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  ram_182 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  ram_183 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  ram_184 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  ram_185 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  ram_186 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  ram_187 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  ram_188 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  ram_189 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  ram_190 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  ram_191 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  ram_192 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  ram_193 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  ram_194 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  ram_195 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  ram_196 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  ram_197 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  ram_198 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  ram_199 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  ram_200 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  ram_201 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  ram_202 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  ram_203 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  ram_204 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  ram_205 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  ram_206 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  ram_207 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  ram_208 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  ram_209 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  ram_210 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  ram_211 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  ram_212 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  ram_213 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  ram_214 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  ram_215 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  ram_216 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  ram_217 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  ram_218 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  ram_219 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  ram_220 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  ram_221 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  ram_222 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  ram_223 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  ram_224 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  ram_225 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  ram_226 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  ram_227 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  ram_228 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  ram_229 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  ram_230 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  ram_231 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  ram_232 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  ram_233 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  ram_234 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  ram_235 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  ram_236 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  ram_237 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  ram_238 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  ram_239 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  ram_240 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  ram_241 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  ram_242 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  ram_243 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  ram_244 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  ram_245 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  ram_246 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  ram_247 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  ram_248 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  ram_249 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  ram_250 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  ram_251 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  ram_252 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  ram_253 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  ram_254 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  ram_255 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  ram_256 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  ram_257 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  ram_258 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  ram_259 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  ram_260 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  ram_261 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  ram_262 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  ram_263 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  ram_264 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  ram_265 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  ram_266 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  ram_267 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  ram_268 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  ram_269 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  ram_270 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  ram_271 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  ram_272 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  ram_273 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  ram_274 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  ram_275 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  ram_276 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  ram_277 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  ram_278 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  ram_279 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  ram_280 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  ram_281 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  ram_282 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  ram_283 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  ram_284 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  ram_285 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  ram_286 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  ram_287 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  ram_288 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  ram_289 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  ram_290 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  ram_291 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  ram_292 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  ram_293 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  ram_294 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  ram_295 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  ram_296 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  ram_297 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  ram_298 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  ram_299 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  ram_300 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  ram_301 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  ram_302 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  ram_303 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  ram_304 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  ram_305 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  ram_306 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  ram_307 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  ram_308 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  ram_309 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  ram_310 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  ram_311 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  ram_312 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  ram_313 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  ram_314 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  ram_315 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  ram_316 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  ram_317 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  ram_318 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  ram_319 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  ram_320 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  ram_321 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  ram_322 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  ram_323 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  ram_324 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  ram_325 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  ram_326 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  ram_327 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  ram_328 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  ram_329 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  ram_330 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  ram_331 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  ram_332 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  ram_333 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  ram_334 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  ram_335 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  ram_336 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  ram_337 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  ram_338 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  ram_339 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  ram_340 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  ram_341 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  ram_342 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  ram_343 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  ram_344 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  ram_345 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  ram_346 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  ram_347 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  ram_348 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  ram_349 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  ram_350 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  ram_351 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  ram_352 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  ram_353 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  ram_354 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  ram_355 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  ram_356 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  ram_357 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  ram_358 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  ram_359 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  ram_360 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  ram_361 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  ram_362 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  ram_363 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  ram_364 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  ram_365 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  ram_366 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  ram_367 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  ram_368 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  ram_369 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  ram_370 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  ram_371 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  ram_372 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  ram_373 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  ram_374 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  ram_375 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  ram_376 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  ram_377 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  ram_378 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  ram_379 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  ram_380 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  ram_381 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  ram_382 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  ram_383 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  ram_384 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  ram_385 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  ram_386 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  ram_387 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  ram_388 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  ram_389 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  ram_390 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  ram_391 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  ram_392 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  ram_393 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  ram_394 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  ram_395 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  ram_396 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  ram_397 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  ram_398 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  ram_399 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  ram_400 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  ram_401 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  ram_402 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  ram_403 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  ram_404 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  ram_405 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  ram_406 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  ram_407 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  ram_408 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  ram_409 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  ram_410 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  ram_411 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  ram_412 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  ram_413 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  ram_414 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  ram_415 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  ram_416 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  ram_417 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  ram_418 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  ram_419 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  ram_420 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  ram_421 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  ram_422 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  ram_423 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  ram_424 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  ram_425 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  ram_426 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  ram_427 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  ram_428 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  ram_429 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  ram_430 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  ram_431 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  ram_432 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  ram_433 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  ram_434 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  ram_435 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  ram_436 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  ram_437 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  ram_438 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  ram_439 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  ram_440 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  ram_441 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  ram_442 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  ram_443 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  ram_444 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  ram_445 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  ram_446 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  ram_447 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  ram_448 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  ram_449 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  ram_450 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  ram_451 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  ram_452 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  ram_453 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  ram_454 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  ram_455 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  ram_456 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  ram_457 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  ram_458 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  ram_459 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  ram_460 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  ram_461 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  ram_462 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  ram_463 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  ram_464 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  ram_465 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  ram_466 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  ram_467 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  ram_468 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  ram_469 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  ram_470 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  ram_471 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  ram_472 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  ram_473 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  ram_474 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  ram_475 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  ram_476 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  ram_477 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  ram_478 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  ram_479 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  ram_480 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  ram_481 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  ram_482 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  ram_483 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  ram_484 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  ram_485 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  ram_486 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  ram_487 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  ram_488 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  ram_489 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  ram_490 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  ram_491 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  ram_492 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  ram_493 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  ram_494 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  ram_495 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  ram_496 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  ram_497 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  ram_498 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  ram_499 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  ram_500 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  ram_501 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  ram_502 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  ram_503 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  ram_504 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  ram_505 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  ram_506 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  ram_507 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  ram_508 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  ram_509 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  ram_510 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  ram_511 = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  ram_512 = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  ram_513 = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  ram_514 = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  ram_515 = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  ram_516 = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  ram_517 = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  ram_518 = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  ram_519 = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  ram_520 = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  ram_521 = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  ram_522 = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  ram_523 = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  ram_524 = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  ram_525 = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  ram_526 = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  ram_527 = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  ram_528 = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  ram_529 = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  ram_530 = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  ram_531 = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  ram_532 = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  ram_533 = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  ram_534 = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  ram_535 = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  ram_536 = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  ram_537 = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  ram_538 = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  ram_539 = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  ram_540 = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  ram_541 = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  ram_542 = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  ram_543 = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  ram_544 = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  ram_545 = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  ram_546 = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  ram_547 = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  ram_548 = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  ram_549 = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  ram_550 = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  ram_551 = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  ram_552 = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  ram_553 = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  ram_554 = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  ram_555 = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  ram_556 = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  ram_557 = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  ram_558 = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  ram_559 = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  ram_560 = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  ram_561 = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  ram_562 = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  ram_563 = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  ram_564 = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  ram_565 = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  ram_566 = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  ram_567 = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  ram_568 = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  ram_569 = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  ram_570 = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  ram_571 = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  ram_572 = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  ram_573 = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  ram_574 = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  ram_575 = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  ram_576 = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  ram_577 = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  ram_578 = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  ram_579 = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  ram_580 = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  ram_581 = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  ram_582 = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  ram_583 = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  ram_584 = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  ram_585 = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  ram_586 = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  ram_587 = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  ram_588 = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  ram_589 = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  ram_590 = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  ram_591 = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  ram_592 = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  ram_593 = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  ram_594 = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  ram_595 = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  ram_596 = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  ram_597 = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  ram_598 = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  ram_599 = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  ram_600 = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  ram_601 = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  ram_602 = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  ram_603 = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  ram_604 = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  ram_605 = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  ram_606 = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  ram_607 = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  ram_608 = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  ram_609 = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  ram_610 = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  ram_611 = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  ram_612 = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  ram_613 = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  ram_614 = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  ram_615 = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  ram_616 = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  ram_617 = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  ram_618 = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  ram_619 = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  ram_620 = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  ram_621 = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  ram_622 = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  ram_623 = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  ram_624 = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  ram_625 = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  ram_626 = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  ram_627 = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  ram_628 = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  ram_629 = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  ram_630 = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  ram_631 = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  ram_632 = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  ram_633 = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  ram_634 = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  ram_635 = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  ram_636 = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  ram_637 = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  ram_638 = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  ram_639 = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  ram_640 = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  ram_641 = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  ram_642 = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  ram_643 = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  ram_644 = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  ram_645 = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  ram_646 = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  ram_647 = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  ram_648 = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  ram_649 = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  ram_650 = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  ram_651 = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  ram_652 = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  ram_653 = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  ram_654 = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  ram_655 = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  ram_656 = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  ram_657 = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  ram_658 = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  ram_659 = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  ram_660 = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  ram_661 = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  ram_662 = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  ram_663 = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  ram_664 = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  ram_665 = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  ram_666 = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  ram_667 = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  ram_668 = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  ram_669 = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  ram_670 = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  ram_671 = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  ram_672 = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  ram_673 = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  ram_674 = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  ram_675 = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  ram_676 = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  ram_677 = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  ram_678 = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  ram_679 = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  ram_680 = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  ram_681 = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  ram_682 = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  ram_683 = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  ram_684 = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  ram_685 = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  ram_686 = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  ram_687 = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  ram_688 = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  ram_689 = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  ram_690 = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  ram_691 = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  ram_692 = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  ram_693 = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  ram_694 = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  ram_695 = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  ram_696 = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  ram_697 = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  ram_698 = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  ram_699 = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  ram_700 = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  ram_701 = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  ram_702 = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  ram_703 = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  ram_704 = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  ram_705 = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  ram_706 = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  ram_707 = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  ram_708 = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  ram_709 = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  ram_710 = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  ram_711 = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  ram_712 = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  ram_713 = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  ram_714 = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  ram_715 = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  ram_716 = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  ram_717 = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  ram_718 = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  ram_719 = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  ram_720 = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  ram_721 = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  ram_722 = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  ram_723 = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  ram_724 = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  ram_725 = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  ram_726 = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  ram_727 = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  ram_728 = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  ram_729 = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  ram_730 = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  ram_731 = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  ram_732 = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  ram_733 = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  ram_734 = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  ram_735 = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  ram_736 = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  ram_737 = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  ram_738 = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  ram_739 = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  ram_740 = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  ram_741 = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  ram_742 = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  ram_743 = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  ram_744 = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  ram_745 = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  ram_746 = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  ram_747 = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  ram_748 = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  ram_749 = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  ram_750 = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  ram_751 = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  ram_752 = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  ram_753 = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  ram_754 = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  ram_755 = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  ram_756 = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  ram_757 = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  ram_758 = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  ram_759 = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  ram_760 = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  ram_761 = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  ram_762 = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  ram_763 = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  ram_764 = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  ram_765 = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  ram_766 = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  ram_767 = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  ram_768 = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  ram_769 = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  ram_770 = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  ram_771 = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  ram_772 = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  ram_773 = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  ram_774 = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  ram_775 = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  ram_776 = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  ram_777 = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  ram_778 = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  ram_779 = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  ram_780 = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  ram_781 = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  ram_782 = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  ram_783 = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  ram_784 = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  ram_785 = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  ram_786 = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  ram_787 = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  ram_788 = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  ram_789 = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  ram_790 = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  ram_791 = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  ram_792 = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  ram_793 = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  ram_794 = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  ram_795 = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  ram_796 = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  ram_797 = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  ram_798 = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  ram_799 = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  ram_800 = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  ram_801 = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  ram_802 = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  ram_803 = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  ram_804 = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  ram_805 = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  ram_806 = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  ram_807 = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  ram_808 = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  ram_809 = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  ram_810 = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  ram_811 = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  ram_812 = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  ram_813 = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  ram_814 = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  ram_815 = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  ram_816 = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  ram_817 = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  ram_818 = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  ram_819 = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  ram_820 = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  ram_821 = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  ram_822 = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  ram_823 = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  ram_824 = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  ram_825 = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  ram_826 = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  ram_827 = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  ram_828 = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  ram_829 = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  ram_830 = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  ram_831 = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  ram_832 = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  ram_833 = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  ram_834 = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  ram_835 = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  ram_836 = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  ram_837 = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  ram_838 = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  ram_839 = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  ram_840 = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  ram_841 = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  ram_842 = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  ram_843 = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  ram_844 = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  ram_845 = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  ram_846 = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  ram_847 = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  ram_848 = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  ram_849 = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  ram_850 = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  ram_851 = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  ram_852 = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  ram_853 = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  ram_854 = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  ram_855 = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  ram_856 = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  ram_857 = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  ram_858 = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  ram_859 = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  ram_860 = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  ram_861 = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  ram_862 = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  ram_863 = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  ram_864 = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  ram_865 = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  ram_866 = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  ram_867 = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  ram_868 = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  ram_869 = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  ram_870 = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  ram_871 = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  ram_872 = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  ram_873 = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  ram_874 = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  ram_875 = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  ram_876 = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  ram_877 = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  ram_878 = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  ram_879 = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  ram_880 = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  ram_881 = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  ram_882 = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  ram_883 = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  ram_884 = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  ram_885 = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  ram_886 = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  ram_887 = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  ram_888 = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  ram_889 = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  ram_890 = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  ram_891 = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  ram_892 = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  ram_893 = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  ram_894 = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  ram_895 = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  ram_896 = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  ram_897 = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  ram_898 = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  ram_899 = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  ram_900 = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  ram_901 = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  ram_902 = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  ram_903 = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  ram_904 = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  ram_905 = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  ram_906 = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  ram_907 = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  ram_908 = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  ram_909 = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  ram_910 = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  ram_911 = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  ram_912 = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  ram_913 = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  ram_914 = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  ram_915 = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  ram_916 = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  ram_917 = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  ram_918 = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  ram_919 = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  ram_920 = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  ram_921 = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  ram_922 = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  ram_923 = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  ram_924 = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  ram_925 = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  ram_926 = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  ram_927 = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  ram_928 = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  ram_929 = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  ram_930 = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  ram_931 = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  ram_932 = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  ram_933 = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  ram_934 = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  ram_935 = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  ram_936 = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  ram_937 = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  ram_938 = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  ram_939 = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  ram_940 = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  ram_941 = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  ram_942 = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  ram_943 = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  ram_944 = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  ram_945 = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  ram_946 = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  ram_947 = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  ram_948 = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  ram_949 = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  ram_950 = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  ram_951 = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  ram_952 = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  ram_953 = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  ram_954 = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  ram_955 = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  ram_956 = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  ram_957 = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  ram_958 = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  ram_959 = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  ram_960 = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  ram_961 = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  ram_962 = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  ram_963 = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  ram_964 = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  ram_965 = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  ram_966 = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  ram_967 = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  ram_968 = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  ram_969 = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  ram_970 = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  ram_971 = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  ram_972 = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  ram_973 = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  ram_974 = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  ram_975 = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  ram_976 = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  ram_977 = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  ram_978 = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  ram_979 = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  ram_980 = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  ram_981 = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  ram_982 = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  ram_983 = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  ram_984 = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  ram_985 = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  ram_986 = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  ram_987 = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  ram_988 = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  ram_989 = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  ram_990 = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  ram_991 = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  ram_992 = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  ram_993 = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  ram_994 = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  ram_995 = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  ram_996 = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  ram_997 = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  ram_998 = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  ram_999 = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  ram_1000 = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  ram_1001 = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  ram_1002 = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  ram_1003 = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  ram_1004 = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  ram_1005 = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  ram_1006 = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  ram_1007 = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  ram_1008 = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  ram_1009 = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  ram_1010 = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  ram_1011 = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  ram_1012 = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  ram_1013 = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  ram_1014 = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  ram_1015 = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  ram_1016 = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  ram_1017 = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  ram_1018 = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  ram_1019 = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  ram_1020 = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  ram_1021 = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  ram_1022 = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  ram_1023 = _RAND_1023[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [7:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [7:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:63]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [5:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [7:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [7:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [5:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [5:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [5:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [5:0] _value_T_1 = enq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  wire [5:0] _value_T_3 = deq_ptr_value + 6'h1; // @[Counter.scala 78:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 6'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ParallelInSerialOut(
  input        clock,
  input        reset,
  input  [7:0] io_shiftIn,
  input        io_load,
  input        io_enable,
  output       io_shiftOut
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] reg_; // @[ShiftReg.scala 47:20]
  wire [7:0] _reg_T_1 = {reg_[6:0],1'h1}; // @[Cat.scala 31:58]
  assign io_shiftOut = reg_[7]; // @[ShiftReg.scala 54:21]
  always @(posedge clock) begin
    if (reset) begin // @[ShiftReg.scala 47:20]
      reg_ <= 8'h0; // @[ShiftReg.scala 47:20]
    end else if (io_load) begin // @[ShiftReg.scala 48:17]
      reg_ <= io_shiftIn; // @[ShiftReg.scala 49:9]
    end else if (io_enable) begin // @[ShiftReg.scala 50:25]
      reg_ <= _reg_T_1; // @[ShiftReg.scala 51:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_ = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module UartTx(
  input        clock,
  input        reset,
  output       io_sendData_ready,
  input        io_sendData_valid,
  input  [7:0] io_sendData_bits,
  output       io_txData
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  shiftReg_clock; // @[Uart.scala 87:24]
  wire  shiftReg_reset; // @[Uart.scala 87:24]
  wire [7:0] shiftReg_io_shiftIn; // @[Uart.scala 87:24]
  wire  shiftReg_io_load; // @[Uart.scala 87:24]
  wire  shiftReg_io_enable; // @[Uart.scala 87:24]
  wire  shiftReg_io_shiftOut; // @[Uart.scala 87:24]
  reg [1:0] state; // @[Uart.scala 78:22]
  reg [9:0] txCount; // @[Counter.scala 62:40]
  wire  wrap_wrap = txCount == 10'h25e; // @[Counter.scala 74:24]
  wire [9:0] _wrap_value_T_1 = txCount + 10'h1; // @[Counter.scala 78:24]
  reg [2:0] sendCount; // @[Uart.scala 84:22]
  wire [7:0] _GEN_15 = {{4'd0}, io_sendData_bits[7:4]}; // @[Bitwise.scala 105:31]
  wire [7:0] _shiftReg_io_shiftIn_T_3 = _GEN_15 & 8'hf; // @[Bitwise.scala 105:31]
  wire [7:0] _shiftReg_io_shiftIn_T_5 = {io_sendData_bits[3:0], 4'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _shiftReg_io_shiftIn_T_7 = _shiftReg_io_shiftIn_T_5 & 8'hf0; // @[Bitwise.scala 105:80]
  wire [7:0] _shiftReg_io_shiftIn_T_8 = _shiftReg_io_shiftIn_T_3 | _shiftReg_io_shiftIn_T_7; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_16 = {{2'd0}, _shiftReg_io_shiftIn_T_8[7:2]}; // @[Bitwise.scala 105:31]
  wire [7:0] _shiftReg_io_shiftIn_T_13 = _GEN_16 & 8'h33; // @[Bitwise.scala 105:31]
  wire [7:0] _shiftReg_io_shiftIn_T_15 = {_shiftReg_io_shiftIn_T_8[5:0], 2'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _shiftReg_io_shiftIn_T_17 = _shiftReg_io_shiftIn_T_15 & 8'hcc; // @[Bitwise.scala 105:80]
  wire [7:0] _shiftReg_io_shiftIn_T_18 = _shiftReg_io_shiftIn_T_13 | _shiftReg_io_shiftIn_T_17; // @[Bitwise.scala 105:39]
  wire [7:0] _GEN_17 = {{1'd0}, _shiftReg_io_shiftIn_T_18[7:1]}; // @[Bitwise.scala 105:31]
  wire [7:0] _shiftReg_io_shiftIn_T_23 = _GEN_17 & 8'h55; // @[Bitwise.scala 105:31]
  wire [7:0] _shiftReg_io_shiftIn_T_25 = {_shiftReg_io_shiftIn_T_18[6:0], 1'h0}; // @[Bitwise.scala 105:70]
  wire [7:0] _shiftReg_io_shiftIn_T_27 = _shiftReg_io_shiftIn_T_25 & 8'haa; // @[Bitwise.scala 105:80]
  wire  _shiftReg_io_load_T_1 = state == 2'h0 & io_sendData_valid; // @[Uart.scala 89:39]
  wire  _shiftReg_io_enable_T = state == 2'h2; // @[Uart.scala 90:31]
  wire [2:0] _sendCount_T_1 = sendCount + 3'h1; // @[Uart.scala 110:34]
  wire [1:0] _GEN_3 = sendCount == 3'h7 ? 2'h3 : state; // @[Uart.scala 107:33 108:17 78:22]
  wire [2:0] _GEN_4 = sendCount == 3'h7 ? sendCount : _sendCount_T_1; // @[Uart.scala 107:33 110:21 84:22]
  wire [1:0] _GEN_5 = 2'h3 == state ? 2'h0 : state; // @[Uart.scala 115:15 99:19 78:22]
  wire [1:0] _GEN_6 = 2'h2 == state ? _GEN_3 : _GEN_5; // @[Uart.scala 99:19]
  wire  _io_txData_T = state == 2'h1; // @[Uart.scala 127:14]
  wire  _io_txData_T_4 = _shiftReg_io_enable_T ? shiftReg_io_shiftOut : 1'h1; // @[Mux.scala 101:16]
  ParallelInSerialOut shiftReg ( // @[Uart.scala 87:24]
    .clock(shiftReg_clock),
    .reset(shiftReg_reset),
    .io_shiftIn(shiftReg_io_shiftIn),
    .io_load(shiftReg_io_load),
    .io_enable(shiftReg_io_enable),
    .io_shiftOut(shiftReg_io_shiftOut)
  );
  assign io_sendData_ready = state == 2'h0; // @[Uart.scala 121:30]
  assign io_txData = _io_txData_T ? 1'h0 : _io_txData_T_4; // @[Mux.scala 101:16]
  assign shiftReg_clock = clock;
  assign shiftReg_reset = reset;
  assign shiftReg_io_shiftIn = _shiftReg_io_shiftIn_T_23 | _shiftReg_io_shiftIn_T_27; // @[Bitwise.scala 105:39]
  assign shiftReg_io_load = state == 2'h0 & io_sendData_valid; // @[Uart.scala 89:39]
  assign shiftReg_io_enable = state == 2'h2 & wrap_wrap; // @[Uart.scala 90:41]
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 78:22]
      state <= 2'h0; // @[Uart.scala 78:22]
    end else if (_shiftReg_io_load_T_1) begin // @[Uart.scala 95:46]
      state <= 2'h1; // @[Uart.scala 96:11]
    end else if (wrap_wrap) begin // @[Uart.scala 98:24]
      if (2'h1 == state) begin // @[Uart.scala 99:19]
        state <= 2'h2; // @[Uart.scala 102:15]
      end else begin
        state <= _GEN_6;
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      txCount <= 10'h0; // @[Counter.scala 62:40]
    end else if (_shiftReg_io_load_T_1) begin // @[Uart.scala 95:46]
      txCount <= 10'h0; // @[Uart.scala 97:13]
    end else if (wrap_wrap) begin // @[Counter.scala 88:20]
      txCount <= 10'h0; // @[Counter.scala 88:28]
    end else begin
      txCount <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
    if (!(_shiftReg_io_load_T_1)) begin // @[Uart.scala 95:46]
      if (wrap_wrap) begin // @[Uart.scala 98:24]
        if (2'h1 == state) begin // @[Uart.scala 99:19]
          sendCount <= 3'h0; // @[Uart.scala 103:19]
        end else if (2'h2 == state) begin // @[Uart.scala 99:19]
          sendCount <= _GEN_4;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  txCount = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  sendCount = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Uart(
  input        clock,
  input        reset,
  output       io_txData,
  input        io_sendData_valid,
  input  [7:0] io_sendData_bits
);
  wire  txQueue_clock; // @[Uart.scala 50:23]
  wire  txQueue_reset; // @[Uart.scala 50:23]
  wire  txQueue_io_enq_ready; // @[Uart.scala 50:23]
  wire  txQueue_io_enq_valid; // @[Uart.scala 50:23]
  wire [7:0] txQueue_io_enq_bits; // @[Uart.scala 50:23]
  wire  txQueue_io_deq_ready; // @[Uart.scala 50:23]
  wire  txQueue_io_deq_valid; // @[Uart.scala 50:23]
  wire [7:0] txQueue_io_deq_bits; // @[Uart.scala 50:23]
  wire  uartTx_clock; // @[Uart.scala 54:22]
  wire  uartTx_reset; // @[Uart.scala 54:22]
  wire  uartTx_io_sendData_ready; // @[Uart.scala 54:22]
  wire  uartTx_io_sendData_valid; // @[Uart.scala 54:22]
  wire [7:0] uartTx_io_sendData_bits; // @[Uart.scala 54:22]
  wire  uartTx_io_txData; // @[Uart.scala 54:22]
  Queue txQueue ( // @[Uart.scala 50:23]
    .clock(txQueue_clock),
    .reset(txQueue_reset),
    .io_enq_ready(txQueue_io_enq_ready),
    .io_enq_valid(txQueue_io_enq_valid),
    .io_enq_bits(txQueue_io_enq_bits),
    .io_deq_ready(txQueue_io_deq_ready),
    .io_deq_valid(txQueue_io_deq_valid),
    .io_deq_bits(txQueue_io_deq_bits)
  );
  UartTx uartTx ( // @[Uart.scala 54:22]
    .clock(uartTx_clock),
    .reset(uartTx_reset),
    .io_sendData_ready(uartTx_io_sendData_ready),
    .io_sendData_valid(uartTx_io_sendData_valid),
    .io_sendData_bits(uartTx_io_sendData_bits),
    .io_txData(uartTx_io_txData)
  );
  assign io_txData = uartTx_io_txData; // @[Uart.scala 55:13]
  assign txQueue_clock = clock;
  assign txQueue_reset = reset;
  assign txQueue_io_enq_valid = io_sendData_valid; // @[Uart.scala 51:18]
  assign txQueue_io_enq_bits = io_sendData_bits; // @[Uart.scala 51:18]
  assign txQueue_io_deq_ready = uartTx_io_sendData_ready; // @[Uart.scala 56:22]
  assign uartTx_clock = clock;
  assign uartTx_reset = reset;
  assign uartTx_io_sendData_valid = txQueue_io_deq_valid; // @[Uart.scala 56:22]
  assign uartTx_io_sendData_bits = txQueue_io_deq_bits; // @[Uart.scala 56:22]
endmodule
module Top(
  input   clock,
  input   reset,
  input   io_rxData,
  output  io_txData
);
  wire  slowClock_clk_original; // @[Top.scala 144:25]
  wire  slowClock_clk_new; // @[Top.scala 144:25]
  wire  cpu_clock; // @[Top.scala 151:21]
  wire  cpu_reset; // @[Top.scala 151:21]
  wire [31:0] cpu_io_iData_addr; // @[Top.scala 151:21]
  wire [31:0] cpu_io_iData_inst; // @[Top.scala 151:21]
  wire [31:0] cpu_io_dData_addr; // @[Top.scala 151:21]
  wire [31:0] cpu_io_dData_writeData; // @[Top.scala 151:21]
  wire  cpu_io_dData_writeEnable; // @[Top.scala 151:21]
  wire [31:0] cpu_io_dData_readData; // @[Top.scala 151:21]
  wire [31:0] iData_io_addr; // @[Top.scala 153:23]
  wire [31:0] iData_io_inst; // @[Top.scala 153:23]
  wire  dData_clock; // @[Top.scala 157:23]
  wire  dData_reset; // @[Top.scala 157:23]
  wire [31:0] dData_io_addr; // @[Top.scala 157:23]
  wire [31:0] dData_io_writeData; // @[Top.scala 157:23]
  wire  dData_io_writeEnable; // @[Top.scala 157:23]
  wire [31:0] dData_io_readData; // @[Top.scala 157:23]
  wire  uart_clock; // @[Top.scala 174:22]
  wire  uart_reset; // @[Top.scala 174:22]
  wire  uart_io_txData; // @[Top.scala 174:22]
  wire  uart_io_sendData_valid; // @[Top.scala 174:22]
  wire [7:0] uart_io_sendData_bits; // @[Top.scala 174:22]
  wire  _T_2 = 32'h80001000 <= cpu_io_dData_addr & cpu_io_dData_addr < 32'h80002000; // @[Top.scala 159:42]
  wire  _T_3 = 32'h10000000 == cpu_io_dData_addr; // @[Top.scala 181:24]
  wire [31:0] _GEN_4 = 32'h10000000 == cpu_io_dData_addr ? cpu_io_dData_writeData : 32'h0; // @[Top.scala 181:47 182:29 185:29]
  wire [31:0] _GEN_6 = _T_2 ? dData_io_readData : 32'h0; // @[Top.scala 195:7 196:29 198:29]
  SlowClock slowClock ( // @[Top.scala 144:25]
    .clk_original(slowClock_clk_original),
    .clk_new(slowClock_clk_new)
  );
  RISCV cpu ( // @[Top.scala 151:21]
    .clock(cpu_clock),
    .reset(cpu_reset),
    .io_iData_addr(cpu_io_iData_addr),
    .io_iData_inst(cpu_io_iData_inst),
    .io_dData_addr(cpu_io_dData_addr),
    .io_dData_writeData(cpu_io_dData_writeData),
    .io_dData_writeEnable(cpu_io_dData_writeEnable),
    .io_dData_readData(cpu_io_dData_readData)
  );
  IData iData ( // @[Top.scala 153:23]
    .io_addr(iData_io_addr),
    .io_inst(iData_io_inst)
  );
  DData dData ( // @[Top.scala 157:23]
    .clock(dData_clock),
    .reset(dData_reset),
    .io_addr(dData_io_addr),
    .io_writeData(dData_io_writeData),
    .io_writeEnable(dData_io_writeEnable),
    .io_readData(dData_io_readData)
  );
  Uart uart ( // @[Top.scala 174:22]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_txData(uart_io_txData),
    .io_sendData_valid(uart_io_sendData_valid),
    .io_sendData_bits(uart_io_sendData_bits)
  );
  assign io_txData = uart_io_txData; // @[Top.scala 178:15]
  assign slowClock_clk_original = clock; // @[Top.scala 145:29]
  assign cpu_clock = slowClock_clk_new;
  assign cpu_reset = reset;
  assign cpu_io_iData_inst = iData_io_inst; // @[Top.scala 154:14]
  assign cpu_io_dData_readData = _T_3 ? 32'h0 : _GEN_6; // @[Top.scala 191:47 192:29]
  assign iData_io_addr = cpu_io_iData_addr; // @[Top.scala 154:14]
  assign dData_clock = slowClock_clk_new;
  assign dData_reset = reset;
  assign dData_io_addr = _T_2 ? cpu_io_dData_addr : 32'h0; // @[Top.scala 160:7 161:21 166:21]
  assign dData_io_writeData = _T_2 ? cpu_io_dData_writeData : 32'h0; // @[Top.scala 160:7 163:26 168:26]
  assign dData_io_writeEnable = _T_2 & cpu_io_dData_writeEnable; // @[Top.scala 160:7 164:28 169:28]
  assign uart_clock = slowClock_clk_new;
  assign uart_reset = reset;
  assign uart_io_sendData_valid = 32'h10000000 == cpu_io_dData_addr & cpu_io_dData_writeEnable; // @[Top.scala 181:47 183:30 186:30]
  assign uart_io_sendData_bits = _GEN_4[7:0];
endmodule
